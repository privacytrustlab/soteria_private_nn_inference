
`include "maxpool1.sv"
`include "fc1.sv"
`include "fc2.sv"
`include "dotproduct5.sv"
`include "dotproduct15.sv"


module mlnn
#(
    parameter INPUTSIZE = 784
)
(
    clk,
    rst,
    g_input,
    e_input,
    o
); 

input clk;
input rst;
input bit [INPUTSIZE-1:0] g_input;
input bit [943:0] e_input;
output bit [9:0] o;

bit [675:0] conv1_0_0;
bit [675:0] conv1_res;
bit [168:0] mp1_0;
bit [168:0] mp1_res;
bit [80:0] conv2_0_0;
bit [80:0] conv2_res;
bit [9:0] fc1_res;
bit [9:0] fc2_res;


    dotproduct5 operation_conv0(.clk (clk), .rst (rst), .g_input ({g_input[0], g_input[1], g_input[28], g_input[30], g_input[56]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[0]));
    dotproduct5 operation_conv1(.clk (clk), .rst (rst), .g_input ({g_input[1], g_input[2], g_input[29], g_input[31], g_input[57]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[1]));
    dotproduct5 operation_conv2(.clk (clk), .rst (rst), .g_input ({g_input[2], g_input[3], g_input[30], g_input[32], g_input[58]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[2]));
    dotproduct5 operation_conv3(.clk (clk), .rst (rst), .g_input ({g_input[3], g_input[4], g_input[31], g_input[33], g_input[59]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[3]));
    dotproduct5 operation_conv4(.clk (clk), .rst (rst), .g_input ({g_input[4], g_input[5], g_input[32], g_input[34], g_input[60]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[4]));
    dotproduct5 operation_conv5(.clk (clk), .rst (rst), .g_input ({g_input[5], g_input[6], g_input[33], g_input[35], g_input[61]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[5]));
    dotproduct5 operation_conv6(.clk (clk), .rst (rst), .g_input ({g_input[6], g_input[7], g_input[34], g_input[36], g_input[62]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[6]));
    dotproduct5 operation_conv7(.clk (clk), .rst (rst), .g_input ({g_input[7], g_input[8], g_input[35], g_input[37], g_input[63]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[7]));
    dotproduct5 operation_conv8(.clk (clk), .rst (rst), .g_input ({g_input[8], g_input[9], g_input[36], g_input[38], g_input[64]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[8]));
    dotproduct5 operation_conv9(.clk (clk), .rst (rst), .g_input ({g_input[9], g_input[10], g_input[37], g_input[39], g_input[65]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[9]));
    dotproduct5 operation_conv10(.clk (clk), .rst (rst), .g_input ({g_input[10], g_input[11], g_input[38], g_input[40], g_input[66]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[10]));
    dotproduct5 operation_conv11(.clk (clk), .rst (rst), .g_input ({g_input[11], g_input[12], g_input[39], g_input[41], g_input[67]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[11]));
    dotproduct5 operation_conv12(.clk (clk), .rst (rst), .g_input ({g_input[12], g_input[13], g_input[40], g_input[42], g_input[68]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[12]));
    dotproduct5 operation_conv13(.clk (clk), .rst (rst), .g_input ({g_input[13], g_input[14], g_input[41], g_input[43], g_input[69]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[13]));
    dotproduct5 operation_conv14(.clk (clk), .rst (rst), .g_input ({g_input[14], g_input[15], g_input[42], g_input[44], g_input[70]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[14]));
    dotproduct5 operation_conv15(.clk (clk), .rst (rst), .g_input ({g_input[15], g_input[16], g_input[43], g_input[45], g_input[71]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[15]));
    dotproduct5 operation_conv16(.clk (clk), .rst (rst), .g_input ({g_input[16], g_input[17], g_input[44], g_input[46], g_input[72]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[16]));
    dotproduct5 operation_conv17(.clk (clk), .rst (rst), .g_input ({g_input[17], g_input[18], g_input[45], g_input[47], g_input[73]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[17]));
    dotproduct5 operation_conv18(.clk (clk), .rst (rst), .g_input ({g_input[18], g_input[19], g_input[46], g_input[48], g_input[74]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[18]));
    dotproduct5 operation_conv19(.clk (clk), .rst (rst), .g_input ({g_input[19], g_input[20], g_input[47], g_input[49], g_input[75]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[19]));
    dotproduct5 operation_conv20(.clk (clk), .rst (rst), .g_input ({g_input[20], g_input[21], g_input[48], g_input[50], g_input[76]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[20]));
    dotproduct5 operation_conv21(.clk (clk), .rst (rst), .g_input ({g_input[21], g_input[22], g_input[49], g_input[51], g_input[77]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[21]));
    dotproduct5 operation_conv22(.clk (clk), .rst (rst), .g_input ({g_input[22], g_input[23], g_input[50], g_input[52], g_input[78]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[22]));
    dotproduct5 operation_conv23(.clk (clk), .rst (rst), .g_input ({g_input[23], g_input[24], g_input[51], g_input[53], g_input[79]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[23]));
    dotproduct5 operation_conv24(.clk (clk), .rst (rst), .g_input ({g_input[24], g_input[25], g_input[52], g_input[54], g_input[80]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[24]));
    dotproduct5 operation_conv25(.clk (clk), .rst (rst), .g_input ({g_input[25], g_input[26], g_input[53], g_input[55], g_input[81]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[25]));
    dotproduct5 operation_conv26(.clk (clk), .rst (rst), .g_input ({g_input[28], g_input[29], g_input[56], g_input[58], g_input[84]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[26]));
    dotproduct5 operation_conv27(.clk (clk), .rst (rst), .g_input ({g_input[29], g_input[30], g_input[57], g_input[59], g_input[85]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[27]));
    dotproduct5 operation_conv28(.clk (clk), .rst (rst), .g_input ({g_input[30], g_input[31], g_input[58], g_input[60], g_input[86]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[28]));
    dotproduct5 operation_conv29(.clk (clk), .rst (rst), .g_input ({g_input[31], g_input[32], g_input[59], g_input[61], g_input[87]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[29]));
    dotproduct5 operation_conv30(.clk (clk), .rst (rst), .g_input ({g_input[32], g_input[33], g_input[60], g_input[62], g_input[88]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[30]));
    dotproduct5 operation_conv31(.clk (clk), .rst (rst), .g_input ({g_input[33], g_input[34], g_input[61], g_input[63], g_input[89]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[31]));
    dotproduct5 operation_conv32(.clk (clk), .rst (rst), .g_input ({g_input[34], g_input[35], g_input[62], g_input[64], g_input[90]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[32]));
    dotproduct5 operation_conv33(.clk (clk), .rst (rst), .g_input ({g_input[35], g_input[36], g_input[63], g_input[65], g_input[91]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[33]));
    dotproduct5 operation_conv34(.clk (clk), .rst (rst), .g_input ({g_input[36], g_input[37], g_input[64], g_input[66], g_input[92]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[34]));
    dotproduct5 operation_conv35(.clk (clk), .rst (rst), .g_input ({g_input[37], g_input[38], g_input[65], g_input[67], g_input[93]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[35]));
    dotproduct5 operation_conv36(.clk (clk), .rst (rst), .g_input ({g_input[38], g_input[39], g_input[66], g_input[68], g_input[94]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[36]));
    dotproduct5 operation_conv37(.clk (clk), .rst (rst), .g_input ({g_input[39], g_input[40], g_input[67], g_input[69], g_input[95]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[37]));
    dotproduct5 operation_conv38(.clk (clk), .rst (rst), .g_input ({g_input[40], g_input[41], g_input[68], g_input[70], g_input[96]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[38]));
    dotproduct5 operation_conv39(.clk (clk), .rst (rst), .g_input ({g_input[41], g_input[42], g_input[69], g_input[71], g_input[97]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[39]));
    dotproduct5 operation_conv40(.clk (clk), .rst (rst), .g_input ({g_input[42], g_input[43], g_input[70], g_input[72], g_input[98]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[40]));
    dotproduct5 operation_conv41(.clk (clk), .rst (rst), .g_input ({g_input[43], g_input[44], g_input[71], g_input[73], g_input[99]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[41]));
    dotproduct5 operation_conv42(.clk (clk), .rst (rst), .g_input ({g_input[44], g_input[45], g_input[72], g_input[74], g_input[100]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[42]));
    dotproduct5 operation_conv43(.clk (clk), .rst (rst), .g_input ({g_input[45], g_input[46], g_input[73], g_input[75], g_input[101]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[43]));
    dotproduct5 operation_conv44(.clk (clk), .rst (rst), .g_input ({g_input[46], g_input[47], g_input[74], g_input[76], g_input[102]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[44]));
    dotproduct5 operation_conv45(.clk (clk), .rst (rst), .g_input ({g_input[47], g_input[48], g_input[75], g_input[77], g_input[103]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[45]));
    dotproduct5 operation_conv46(.clk (clk), .rst (rst), .g_input ({g_input[48], g_input[49], g_input[76], g_input[78], g_input[104]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[46]));
    dotproduct5 operation_conv47(.clk (clk), .rst (rst), .g_input ({g_input[49], g_input[50], g_input[77], g_input[79], g_input[105]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[47]));
    dotproduct5 operation_conv48(.clk (clk), .rst (rst), .g_input ({g_input[50], g_input[51], g_input[78], g_input[80], g_input[106]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[48]));
    dotproduct5 operation_conv49(.clk (clk), .rst (rst), .g_input ({g_input[51], g_input[52], g_input[79], g_input[81], g_input[107]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[49]));
    dotproduct5 operation_conv50(.clk (clk), .rst (rst), .g_input ({g_input[52], g_input[53], g_input[80], g_input[82], g_input[108]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[50]));
    dotproduct5 operation_conv51(.clk (clk), .rst (rst), .g_input ({g_input[53], g_input[54], g_input[81], g_input[83], g_input[109]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[51]));
    dotproduct5 operation_conv52(.clk (clk), .rst (rst), .g_input ({g_input[56], g_input[57], g_input[84], g_input[86], g_input[112]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[52]));
    dotproduct5 operation_conv53(.clk (clk), .rst (rst), .g_input ({g_input[57], g_input[58], g_input[85], g_input[87], g_input[113]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[53]));
    dotproduct5 operation_conv54(.clk (clk), .rst (rst), .g_input ({g_input[58], g_input[59], g_input[86], g_input[88], g_input[114]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[54]));
    dotproduct5 operation_conv55(.clk (clk), .rst (rst), .g_input ({g_input[59], g_input[60], g_input[87], g_input[89], g_input[115]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[55]));
    dotproduct5 operation_conv56(.clk (clk), .rst (rst), .g_input ({g_input[60], g_input[61], g_input[88], g_input[90], g_input[116]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[56]));
    dotproduct5 operation_conv57(.clk (clk), .rst (rst), .g_input ({g_input[61], g_input[62], g_input[89], g_input[91], g_input[117]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[57]));
    dotproduct5 operation_conv58(.clk (clk), .rst (rst), .g_input ({g_input[62], g_input[63], g_input[90], g_input[92], g_input[118]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[58]));
    dotproduct5 operation_conv59(.clk (clk), .rst (rst), .g_input ({g_input[63], g_input[64], g_input[91], g_input[93], g_input[119]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[59]));
    dotproduct5 operation_conv60(.clk (clk), .rst (rst), .g_input ({g_input[64], g_input[65], g_input[92], g_input[94], g_input[120]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[60]));
    dotproduct5 operation_conv61(.clk (clk), .rst (rst), .g_input ({g_input[65], g_input[66], g_input[93], g_input[95], g_input[121]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[61]));
    dotproduct5 operation_conv62(.clk (clk), .rst (rst), .g_input ({g_input[66], g_input[67], g_input[94], g_input[96], g_input[122]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[62]));
    dotproduct5 operation_conv63(.clk (clk), .rst (rst), .g_input ({g_input[67], g_input[68], g_input[95], g_input[97], g_input[123]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[63]));
    dotproduct5 operation_conv64(.clk (clk), .rst (rst), .g_input ({g_input[68], g_input[69], g_input[96], g_input[98], g_input[124]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[64]));
    dotproduct5 operation_conv65(.clk (clk), .rst (rst), .g_input ({g_input[69], g_input[70], g_input[97], g_input[99], g_input[125]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[65]));
    dotproduct5 operation_conv66(.clk (clk), .rst (rst), .g_input ({g_input[70], g_input[71], g_input[98], g_input[100], g_input[126]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[66]));
    dotproduct5 operation_conv67(.clk (clk), .rst (rst), .g_input ({g_input[71], g_input[72], g_input[99], g_input[101], g_input[127]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[67]));
    dotproduct5 operation_conv68(.clk (clk), .rst (rst), .g_input ({g_input[72], g_input[73], g_input[100], g_input[102], g_input[128]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[68]));
    dotproduct5 operation_conv69(.clk (clk), .rst (rst), .g_input ({g_input[73], g_input[74], g_input[101], g_input[103], g_input[129]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[69]));
    dotproduct5 operation_conv70(.clk (clk), .rst (rst), .g_input ({g_input[74], g_input[75], g_input[102], g_input[104], g_input[130]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[70]));
    dotproduct5 operation_conv71(.clk (clk), .rst (rst), .g_input ({g_input[75], g_input[76], g_input[103], g_input[105], g_input[131]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[71]));
    dotproduct5 operation_conv72(.clk (clk), .rst (rst), .g_input ({g_input[76], g_input[77], g_input[104], g_input[106], g_input[132]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[72]));
    dotproduct5 operation_conv73(.clk (clk), .rst (rst), .g_input ({g_input[77], g_input[78], g_input[105], g_input[107], g_input[133]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[73]));
    dotproduct5 operation_conv74(.clk (clk), .rst (rst), .g_input ({g_input[78], g_input[79], g_input[106], g_input[108], g_input[134]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[74]));
    dotproduct5 operation_conv75(.clk (clk), .rst (rst), .g_input ({g_input[79], g_input[80], g_input[107], g_input[109], g_input[135]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[75]));
    dotproduct5 operation_conv76(.clk (clk), .rst (rst), .g_input ({g_input[80], g_input[81], g_input[108], g_input[110], g_input[136]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[76]));
    dotproduct5 operation_conv77(.clk (clk), .rst (rst), .g_input ({g_input[81], g_input[82], g_input[109], g_input[111], g_input[137]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[77]));
    dotproduct5 operation_conv78(.clk (clk), .rst (rst), .g_input ({g_input[84], g_input[85], g_input[112], g_input[114], g_input[140]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[78]));
    dotproduct5 operation_conv79(.clk (clk), .rst (rst), .g_input ({g_input[85], g_input[86], g_input[113], g_input[115], g_input[141]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[79]));
    dotproduct5 operation_conv80(.clk (clk), .rst (rst), .g_input ({g_input[86], g_input[87], g_input[114], g_input[116], g_input[142]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[80]));
    dotproduct5 operation_conv81(.clk (clk), .rst (rst), .g_input ({g_input[87], g_input[88], g_input[115], g_input[117], g_input[143]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[81]));
    dotproduct5 operation_conv82(.clk (clk), .rst (rst), .g_input ({g_input[88], g_input[89], g_input[116], g_input[118], g_input[144]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[82]));
    dotproduct5 operation_conv83(.clk (clk), .rst (rst), .g_input ({g_input[89], g_input[90], g_input[117], g_input[119], g_input[145]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[83]));
    dotproduct5 operation_conv84(.clk (clk), .rst (rst), .g_input ({g_input[90], g_input[91], g_input[118], g_input[120], g_input[146]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[84]));
    dotproduct5 operation_conv85(.clk (clk), .rst (rst), .g_input ({g_input[91], g_input[92], g_input[119], g_input[121], g_input[147]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[85]));
    dotproduct5 operation_conv86(.clk (clk), .rst (rst), .g_input ({g_input[92], g_input[93], g_input[120], g_input[122], g_input[148]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[86]));
    dotproduct5 operation_conv87(.clk (clk), .rst (rst), .g_input ({g_input[93], g_input[94], g_input[121], g_input[123], g_input[149]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[87]));
    dotproduct5 operation_conv88(.clk (clk), .rst (rst), .g_input ({g_input[94], g_input[95], g_input[122], g_input[124], g_input[150]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[88]));
    dotproduct5 operation_conv89(.clk (clk), .rst (rst), .g_input ({g_input[95], g_input[96], g_input[123], g_input[125], g_input[151]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[89]));
    dotproduct5 operation_conv90(.clk (clk), .rst (rst), .g_input ({g_input[96], g_input[97], g_input[124], g_input[126], g_input[152]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[90]));
    dotproduct5 operation_conv91(.clk (clk), .rst (rst), .g_input ({g_input[97], g_input[98], g_input[125], g_input[127], g_input[153]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[91]));
    dotproduct5 operation_conv92(.clk (clk), .rst (rst), .g_input ({g_input[98], g_input[99], g_input[126], g_input[128], g_input[154]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[92]));
    dotproduct5 operation_conv93(.clk (clk), .rst (rst), .g_input ({g_input[99], g_input[100], g_input[127], g_input[129], g_input[155]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[93]));
    dotproduct5 operation_conv94(.clk (clk), .rst (rst), .g_input ({g_input[100], g_input[101], g_input[128], g_input[130], g_input[156]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[94]));
    dotproduct5 operation_conv95(.clk (clk), .rst (rst), .g_input ({g_input[101], g_input[102], g_input[129], g_input[131], g_input[157]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[95]));
    dotproduct5 operation_conv96(.clk (clk), .rst (rst), .g_input ({g_input[102], g_input[103], g_input[130], g_input[132], g_input[158]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[96]));
    dotproduct5 operation_conv97(.clk (clk), .rst (rst), .g_input ({g_input[103], g_input[104], g_input[131], g_input[133], g_input[159]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[97]));
    dotproduct5 operation_conv98(.clk (clk), .rst (rst), .g_input ({g_input[104], g_input[105], g_input[132], g_input[134], g_input[160]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[98]));
    dotproduct5 operation_conv99(.clk (clk), .rst (rst), .g_input ({g_input[105], g_input[106], g_input[133], g_input[135], g_input[161]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[99]));
    dotproduct5 operation_conv100(.clk (clk), .rst (rst), .g_input ({g_input[106], g_input[107], g_input[134], g_input[136], g_input[162]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[100]));
    dotproduct5 operation_conv101(.clk (clk), .rst (rst), .g_input ({g_input[107], g_input[108], g_input[135], g_input[137], g_input[163]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[101]));
    dotproduct5 operation_conv102(.clk (clk), .rst (rst), .g_input ({g_input[108], g_input[109], g_input[136], g_input[138], g_input[164]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[102]));
    dotproduct5 operation_conv103(.clk (clk), .rst (rst), .g_input ({g_input[109], g_input[110], g_input[137], g_input[139], g_input[165]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[103]));
    dotproduct5 operation_conv104(.clk (clk), .rst (rst), .g_input ({g_input[112], g_input[113], g_input[140], g_input[142], g_input[168]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[104]));
    dotproduct5 operation_conv105(.clk (clk), .rst (rst), .g_input ({g_input[113], g_input[114], g_input[141], g_input[143], g_input[169]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[105]));
    dotproduct5 operation_conv106(.clk (clk), .rst (rst), .g_input ({g_input[114], g_input[115], g_input[142], g_input[144], g_input[170]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[106]));
    dotproduct5 operation_conv107(.clk (clk), .rst (rst), .g_input ({g_input[115], g_input[116], g_input[143], g_input[145], g_input[171]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[107]));
    dotproduct5 operation_conv108(.clk (clk), .rst (rst), .g_input ({g_input[116], g_input[117], g_input[144], g_input[146], g_input[172]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[108]));
    dotproduct5 operation_conv109(.clk (clk), .rst (rst), .g_input ({g_input[117], g_input[118], g_input[145], g_input[147], g_input[173]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[109]));
    dotproduct5 operation_conv110(.clk (clk), .rst (rst), .g_input ({g_input[118], g_input[119], g_input[146], g_input[148], g_input[174]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[110]));
    dotproduct5 operation_conv111(.clk (clk), .rst (rst), .g_input ({g_input[119], g_input[120], g_input[147], g_input[149], g_input[175]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[111]));
    dotproduct5 operation_conv112(.clk (clk), .rst (rst), .g_input ({g_input[120], g_input[121], g_input[148], g_input[150], g_input[176]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[112]));
    dotproduct5 operation_conv113(.clk (clk), .rst (rst), .g_input ({g_input[121], g_input[122], g_input[149], g_input[151], g_input[177]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[113]));
    dotproduct5 operation_conv114(.clk (clk), .rst (rst), .g_input ({g_input[122], g_input[123], g_input[150], g_input[152], g_input[178]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[114]));
    dotproduct5 operation_conv115(.clk (clk), .rst (rst), .g_input ({g_input[123], g_input[124], g_input[151], g_input[153], g_input[179]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[115]));
    dotproduct5 operation_conv116(.clk (clk), .rst (rst), .g_input ({g_input[124], g_input[125], g_input[152], g_input[154], g_input[180]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[116]));
    dotproduct5 operation_conv117(.clk (clk), .rst (rst), .g_input ({g_input[125], g_input[126], g_input[153], g_input[155], g_input[181]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[117]));
    dotproduct5 operation_conv118(.clk (clk), .rst (rst), .g_input ({g_input[126], g_input[127], g_input[154], g_input[156], g_input[182]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[118]));
    dotproduct5 operation_conv119(.clk (clk), .rst (rst), .g_input ({g_input[127], g_input[128], g_input[155], g_input[157], g_input[183]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[119]));
    dotproduct5 operation_conv120(.clk (clk), .rst (rst), .g_input ({g_input[128], g_input[129], g_input[156], g_input[158], g_input[184]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[120]));
    dotproduct5 operation_conv121(.clk (clk), .rst (rst), .g_input ({g_input[129], g_input[130], g_input[157], g_input[159], g_input[185]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[121]));
    dotproduct5 operation_conv122(.clk (clk), .rst (rst), .g_input ({g_input[130], g_input[131], g_input[158], g_input[160], g_input[186]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[122]));
    dotproduct5 operation_conv123(.clk (clk), .rst (rst), .g_input ({g_input[131], g_input[132], g_input[159], g_input[161], g_input[187]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[123]));
    dotproduct5 operation_conv124(.clk (clk), .rst (rst), .g_input ({g_input[132], g_input[133], g_input[160], g_input[162], g_input[188]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[124]));
    dotproduct5 operation_conv125(.clk (clk), .rst (rst), .g_input ({g_input[133], g_input[134], g_input[161], g_input[163], g_input[189]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[125]));
    dotproduct5 operation_conv126(.clk (clk), .rst (rst), .g_input ({g_input[134], g_input[135], g_input[162], g_input[164], g_input[190]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[126]));
    dotproduct5 operation_conv127(.clk (clk), .rst (rst), .g_input ({g_input[135], g_input[136], g_input[163], g_input[165], g_input[191]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[127]));
    dotproduct5 operation_conv128(.clk (clk), .rst (rst), .g_input ({g_input[136], g_input[137], g_input[164], g_input[166], g_input[192]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[128]));
    dotproduct5 operation_conv129(.clk (clk), .rst (rst), .g_input ({g_input[137], g_input[138], g_input[165], g_input[167], g_input[193]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[129]));
    dotproduct5 operation_conv130(.clk (clk), .rst (rst), .g_input ({g_input[140], g_input[141], g_input[168], g_input[170], g_input[196]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[130]));
    dotproduct5 operation_conv131(.clk (clk), .rst (rst), .g_input ({g_input[141], g_input[142], g_input[169], g_input[171], g_input[197]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[131]));
    dotproduct5 operation_conv132(.clk (clk), .rst (rst), .g_input ({g_input[142], g_input[143], g_input[170], g_input[172], g_input[198]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[132]));
    dotproduct5 operation_conv133(.clk (clk), .rst (rst), .g_input ({g_input[143], g_input[144], g_input[171], g_input[173], g_input[199]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[133]));
    dotproduct5 operation_conv134(.clk (clk), .rst (rst), .g_input ({g_input[144], g_input[145], g_input[172], g_input[174], g_input[200]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[134]));
    dotproduct5 operation_conv135(.clk (clk), .rst (rst), .g_input ({g_input[145], g_input[146], g_input[173], g_input[175], g_input[201]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[135]));
    dotproduct5 operation_conv136(.clk (clk), .rst (rst), .g_input ({g_input[146], g_input[147], g_input[174], g_input[176], g_input[202]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[136]));
    dotproduct5 operation_conv137(.clk (clk), .rst (rst), .g_input ({g_input[147], g_input[148], g_input[175], g_input[177], g_input[203]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[137]));
    dotproduct5 operation_conv138(.clk (clk), .rst (rst), .g_input ({g_input[148], g_input[149], g_input[176], g_input[178], g_input[204]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[138]));
    dotproduct5 operation_conv139(.clk (clk), .rst (rst), .g_input ({g_input[149], g_input[150], g_input[177], g_input[179], g_input[205]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[139]));
    dotproduct5 operation_conv140(.clk (clk), .rst (rst), .g_input ({g_input[150], g_input[151], g_input[178], g_input[180], g_input[206]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[140]));
    dotproduct5 operation_conv141(.clk (clk), .rst (rst), .g_input ({g_input[151], g_input[152], g_input[179], g_input[181], g_input[207]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[141]));
    dotproduct5 operation_conv142(.clk (clk), .rst (rst), .g_input ({g_input[152], g_input[153], g_input[180], g_input[182], g_input[208]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[142]));
    dotproduct5 operation_conv143(.clk (clk), .rst (rst), .g_input ({g_input[153], g_input[154], g_input[181], g_input[183], g_input[209]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[143]));
    dotproduct5 operation_conv144(.clk (clk), .rst (rst), .g_input ({g_input[154], g_input[155], g_input[182], g_input[184], g_input[210]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[144]));
    dotproduct5 operation_conv145(.clk (clk), .rst (rst), .g_input ({g_input[155], g_input[156], g_input[183], g_input[185], g_input[211]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[145]));
    dotproduct5 operation_conv146(.clk (clk), .rst (rst), .g_input ({g_input[156], g_input[157], g_input[184], g_input[186], g_input[212]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[146]));
    dotproduct5 operation_conv147(.clk (clk), .rst (rst), .g_input ({g_input[157], g_input[158], g_input[185], g_input[187], g_input[213]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[147]));
    dotproduct5 operation_conv148(.clk (clk), .rst (rst), .g_input ({g_input[158], g_input[159], g_input[186], g_input[188], g_input[214]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[148]));
    dotproduct5 operation_conv149(.clk (clk), .rst (rst), .g_input ({g_input[159], g_input[160], g_input[187], g_input[189], g_input[215]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[149]));
    dotproduct5 operation_conv150(.clk (clk), .rst (rst), .g_input ({g_input[160], g_input[161], g_input[188], g_input[190], g_input[216]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[150]));
    dotproduct5 operation_conv151(.clk (clk), .rst (rst), .g_input ({g_input[161], g_input[162], g_input[189], g_input[191], g_input[217]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[151]));
    dotproduct5 operation_conv152(.clk (clk), .rst (rst), .g_input ({g_input[162], g_input[163], g_input[190], g_input[192], g_input[218]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[152]));
    dotproduct5 operation_conv153(.clk (clk), .rst (rst), .g_input ({g_input[163], g_input[164], g_input[191], g_input[193], g_input[219]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[153]));
    dotproduct5 operation_conv154(.clk (clk), .rst (rst), .g_input ({g_input[164], g_input[165], g_input[192], g_input[194], g_input[220]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[154]));
    dotproduct5 operation_conv155(.clk (clk), .rst (rst), .g_input ({g_input[165], g_input[166], g_input[193], g_input[195], g_input[221]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[155]));
    dotproduct5 operation_conv156(.clk (clk), .rst (rst), .g_input ({g_input[168], g_input[169], g_input[196], g_input[198], g_input[224]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[156]));
    dotproduct5 operation_conv157(.clk (clk), .rst (rst), .g_input ({g_input[169], g_input[170], g_input[197], g_input[199], g_input[225]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[157]));
    dotproduct5 operation_conv158(.clk (clk), .rst (rst), .g_input ({g_input[170], g_input[171], g_input[198], g_input[200], g_input[226]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[158]));
    dotproduct5 operation_conv159(.clk (clk), .rst (rst), .g_input ({g_input[171], g_input[172], g_input[199], g_input[201], g_input[227]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[159]));
    dotproduct5 operation_conv160(.clk (clk), .rst (rst), .g_input ({g_input[172], g_input[173], g_input[200], g_input[202], g_input[228]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[160]));
    dotproduct5 operation_conv161(.clk (clk), .rst (rst), .g_input ({g_input[173], g_input[174], g_input[201], g_input[203], g_input[229]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[161]));
    dotproduct5 operation_conv162(.clk (clk), .rst (rst), .g_input ({g_input[174], g_input[175], g_input[202], g_input[204], g_input[230]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[162]));
    dotproduct5 operation_conv163(.clk (clk), .rst (rst), .g_input ({g_input[175], g_input[176], g_input[203], g_input[205], g_input[231]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[163]));
    dotproduct5 operation_conv164(.clk (clk), .rst (rst), .g_input ({g_input[176], g_input[177], g_input[204], g_input[206], g_input[232]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[164]));
    dotproduct5 operation_conv165(.clk (clk), .rst (rst), .g_input ({g_input[177], g_input[178], g_input[205], g_input[207], g_input[233]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[165]));
    dotproduct5 operation_conv166(.clk (clk), .rst (rst), .g_input ({g_input[178], g_input[179], g_input[206], g_input[208], g_input[234]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[166]));
    dotproduct5 operation_conv167(.clk (clk), .rst (rst), .g_input ({g_input[179], g_input[180], g_input[207], g_input[209], g_input[235]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[167]));
    dotproduct5 operation_conv168(.clk (clk), .rst (rst), .g_input ({g_input[180], g_input[181], g_input[208], g_input[210], g_input[236]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[168]));
    dotproduct5 operation_conv169(.clk (clk), .rst (rst), .g_input ({g_input[181], g_input[182], g_input[209], g_input[211], g_input[237]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[169]));
    dotproduct5 operation_conv170(.clk (clk), .rst (rst), .g_input ({g_input[182], g_input[183], g_input[210], g_input[212], g_input[238]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[170]));
    dotproduct5 operation_conv171(.clk (clk), .rst (rst), .g_input ({g_input[183], g_input[184], g_input[211], g_input[213], g_input[239]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[171]));
    dotproduct5 operation_conv172(.clk (clk), .rst (rst), .g_input ({g_input[184], g_input[185], g_input[212], g_input[214], g_input[240]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[172]));
    dotproduct5 operation_conv173(.clk (clk), .rst (rst), .g_input ({g_input[185], g_input[186], g_input[213], g_input[215], g_input[241]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[173]));
    dotproduct5 operation_conv174(.clk (clk), .rst (rst), .g_input ({g_input[186], g_input[187], g_input[214], g_input[216], g_input[242]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[174]));
    dotproduct5 operation_conv175(.clk (clk), .rst (rst), .g_input ({g_input[187], g_input[188], g_input[215], g_input[217], g_input[243]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[175]));
    dotproduct5 operation_conv176(.clk (clk), .rst (rst), .g_input ({g_input[188], g_input[189], g_input[216], g_input[218], g_input[244]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[176]));
    dotproduct5 operation_conv177(.clk (clk), .rst (rst), .g_input ({g_input[189], g_input[190], g_input[217], g_input[219], g_input[245]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[177]));
    dotproduct5 operation_conv178(.clk (clk), .rst (rst), .g_input ({g_input[190], g_input[191], g_input[218], g_input[220], g_input[246]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[178]));
    dotproduct5 operation_conv179(.clk (clk), .rst (rst), .g_input ({g_input[191], g_input[192], g_input[219], g_input[221], g_input[247]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[179]));
    dotproduct5 operation_conv180(.clk (clk), .rst (rst), .g_input ({g_input[192], g_input[193], g_input[220], g_input[222], g_input[248]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[180]));
    dotproduct5 operation_conv181(.clk (clk), .rst (rst), .g_input ({g_input[193], g_input[194], g_input[221], g_input[223], g_input[249]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[181]));
    dotproduct5 operation_conv182(.clk (clk), .rst (rst), .g_input ({g_input[196], g_input[197], g_input[224], g_input[226], g_input[252]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[182]));
    dotproduct5 operation_conv183(.clk (clk), .rst (rst), .g_input ({g_input[197], g_input[198], g_input[225], g_input[227], g_input[253]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[183]));
    dotproduct5 operation_conv184(.clk (clk), .rst (rst), .g_input ({g_input[198], g_input[199], g_input[226], g_input[228], g_input[254]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[184]));
    dotproduct5 operation_conv185(.clk (clk), .rst (rst), .g_input ({g_input[199], g_input[200], g_input[227], g_input[229], g_input[255]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[185]));
    dotproduct5 operation_conv186(.clk (clk), .rst (rst), .g_input ({g_input[200], g_input[201], g_input[228], g_input[230], g_input[256]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[186]));
    dotproduct5 operation_conv187(.clk (clk), .rst (rst), .g_input ({g_input[201], g_input[202], g_input[229], g_input[231], g_input[257]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[187]));
    dotproduct5 operation_conv188(.clk (clk), .rst (rst), .g_input ({g_input[202], g_input[203], g_input[230], g_input[232], g_input[258]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[188]));
    dotproduct5 operation_conv189(.clk (clk), .rst (rst), .g_input ({g_input[203], g_input[204], g_input[231], g_input[233], g_input[259]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[189]));
    dotproduct5 operation_conv190(.clk (clk), .rst (rst), .g_input ({g_input[204], g_input[205], g_input[232], g_input[234], g_input[260]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[190]));
    dotproduct5 operation_conv191(.clk (clk), .rst (rst), .g_input ({g_input[205], g_input[206], g_input[233], g_input[235], g_input[261]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[191]));
    dotproduct5 operation_conv192(.clk (clk), .rst (rst), .g_input ({g_input[206], g_input[207], g_input[234], g_input[236], g_input[262]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[192]));
    dotproduct5 operation_conv193(.clk (clk), .rst (rst), .g_input ({g_input[207], g_input[208], g_input[235], g_input[237], g_input[263]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[193]));
    dotproduct5 operation_conv194(.clk (clk), .rst (rst), .g_input ({g_input[208], g_input[209], g_input[236], g_input[238], g_input[264]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[194]));
    dotproduct5 operation_conv195(.clk (clk), .rst (rst), .g_input ({g_input[209], g_input[210], g_input[237], g_input[239], g_input[265]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[195]));
    dotproduct5 operation_conv196(.clk (clk), .rst (rst), .g_input ({g_input[210], g_input[211], g_input[238], g_input[240], g_input[266]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[196]));
    dotproduct5 operation_conv197(.clk (clk), .rst (rst), .g_input ({g_input[211], g_input[212], g_input[239], g_input[241], g_input[267]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[197]));
    dotproduct5 operation_conv198(.clk (clk), .rst (rst), .g_input ({g_input[212], g_input[213], g_input[240], g_input[242], g_input[268]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[198]));
    dotproduct5 operation_conv199(.clk (clk), .rst (rst), .g_input ({g_input[213], g_input[214], g_input[241], g_input[243], g_input[269]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[199]));
    dotproduct5 operation_conv200(.clk (clk), .rst (rst), .g_input ({g_input[214], g_input[215], g_input[242], g_input[244], g_input[270]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[200]));
    dotproduct5 operation_conv201(.clk (clk), .rst (rst), .g_input ({g_input[215], g_input[216], g_input[243], g_input[245], g_input[271]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[201]));
    dotproduct5 operation_conv202(.clk (clk), .rst (rst), .g_input ({g_input[216], g_input[217], g_input[244], g_input[246], g_input[272]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[202]));
    dotproduct5 operation_conv203(.clk (clk), .rst (rst), .g_input ({g_input[217], g_input[218], g_input[245], g_input[247], g_input[273]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[203]));
    dotproduct5 operation_conv204(.clk (clk), .rst (rst), .g_input ({g_input[218], g_input[219], g_input[246], g_input[248], g_input[274]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[204]));
    dotproduct5 operation_conv205(.clk (clk), .rst (rst), .g_input ({g_input[219], g_input[220], g_input[247], g_input[249], g_input[275]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[205]));
    dotproduct5 operation_conv206(.clk (clk), .rst (rst), .g_input ({g_input[220], g_input[221], g_input[248], g_input[250], g_input[276]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[206]));
    dotproduct5 operation_conv207(.clk (clk), .rst (rst), .g_input ({g_input[221], g_input[222], g_input[249], g_input[251], g_input[277]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[207]));
    dotproduct5 operation_conv208(.clk (clk), .rst (rst), .g_input ({g_input[224], g_input[225], g_input[252], g_input[254], g_input[280]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[208]));
    dotproduct5 operation_conv209(.clk (clk), .rst (rst), .g_input ({g_input[225], g_input[226], g_input[253], g_input[255], g_input[281]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[209]));
    dotproduct5 operation_conv210(.clk (clk), .rst (rst), .g_input ({g_input[226], g_input[227], g_input[254], g_input[256], g_input[282]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[210]));
    dotproduct5 operation_conv211(.clk (clk), .rst (rst), .g_input ({g_input[227], g_input[228], g_input[255], g_input[257], g_input[283]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[211]));
    dotproduct5 operation_conv212(.clk (clk), .rst (rst), .g_input ({g_input[228], g_input[229], g_input[256], g_input[258], g_input[284]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[212]));
    dotproduct5 operation_conv213(.clk (clk), .rst (rst), .g_input ({g_input[229], g_input[230], g_input[257], g_input[259], g_input[285]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[213]));
    dotproduct5 operation_conv214(.clk (clk), .rst (rst), .g_input ({g_input[230], g_input[231], g_input[258], g_input[260], g_input[286]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[214]));
    dotproduct5 operation_conv215(.clk (clk), .rst (rst), .g_input ({g_input[231], g_input[232], g_input[259], g_input[261], g_input[287]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[215]));
    dotproduct5 operation_conv216(.clk (clk), .rst (rst), .g_input ({g_input[232], g_input[233], g_input[260], g_input[262], g_input[288]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[216]));
    dotproduct5 operation_conv217(.clk (clk), .rst (rst), .g_input ({g_input[233], g_input[234], g_input[261], g_input[263], g_input[289]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[217]));
    dotproduct5 operation_conv218(.clk (clk), .rst (rst), .g_input ({g_input[234], g_input[235], g_input[262], g_input[264], g_input[290]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[218]));
    dotproduct5 operation_conv219(.clk (clk), .rst (rst), .g_input ({g_input[235], g_input[236], g_input[263], g_input[265], g_input[291]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[219]));
    dotproduct5 operation_conv220(.clk (clk), .rst (rst), .g_input ({g_input[236], g_input[237], g_input[264], g_input[266], g_input[292]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[220]));
    dotproduct5 operation_conv221(.clk (clk), .rst (rst), .g_input ({g_input[237], g_input[238], g_input[265], g_input[267], g_input[293]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[221]));
    dotproduct5 operation_conv222(.clk (clk), .rst (rst), .g_input ({g_input[238], g_input[239], g_input[266], g_input[268], g_input[294]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[222]));
    dotproduct5 operation_conv223(.clk (clk), .rst (rst), .g_input ({g_input[239], g_input[240], g_input[267], g_input[269], g_input[295]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[223]));
    dotproduct5 operation_conv224(.clk (clk), .rst (rst), .g_input ({g_input[240], g_input[241], g_input[268], g_input[270], g_input[296]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[224]));
    dotproduct5 operation_conv225(.clk (clk), .rst (rst), .g_input ({g_input[241], g_input[242], g_input[269], g_input[271], g_input[297]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[225]));
    dotproduct5 operation_conv226(.clk (clk), .rst (rst), .g_input ({g_input[242], g_input[243], g_input[270], g_input[272], g_input[298]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[226]));
    dotproduct5 operation_conv227(.clk (clk), .rst (rst), .g_input ({g_input[243], g_input[244], g_input[271], g_input[273], g_input[299]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[227]));
    dotproduct5 operation_conv228(.clk (clk), .rst (rst), .g_input ({g_input[244], g_input[245], g_input[272], g_input[274], g_input[300]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[228]));
    dotproduct5 operation_conv229(.clk (clk), .rst (rst), .g_input ({g_input[245], g_input[246], g_input[273], g_input[275], g_input[301]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[229]));
    dotproduct5 operation_conv230(.clk (clk), .rst (rst), .g_input ({g_input[246], g_input[247], g_input[274], g_input[276], g_input[302]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[230]));
    dotproduct5 operation_conv231(.clk (clk), .rst (rst), .g_input ({g_input[247], g_input[248], g_input[275], g_input[277], g_input[303]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[231]));
    dotproduct5 operation_conv232(.clk (clk), .rst (rst), .g_input ({g_input[248], g_input[249], g_input[276], g_input[278], g_input[304]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[232]));
    dotproduct5 operation_conv233(.clk (clk), .rst (rst), .g_input ({g_input[249], g_input[250], g_input[277], g_input[279], g_input[305]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[233]));
    dotproduct5 operation_conv234(.clk (clk), .rst (rst), .g_input ({g_input[252], g_input[253], g_input[280], g_input[282], g_input[308]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[234]));
    dotproduct5 operation_conv235(.clk (clk), .rst (rst), .g_input ({g_input[253], g_input[254], g_input[281], g_input[283], g_input[309]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[235]));
    dotproduct5 operation_conv236(.clk (clk), .rst (rst), .g_input ({g_input[254], g_input[255], g_input[282], g_input[284], g_input[310]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[236]));
    dotproduct5 operation_conv237(.clk (clk), .rst (rst), .g_input ({g_input[255], g_input[256], g_input[283], g_input[285], g_input[311]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[237]));
    dotproduct5 operation_conv238(.clk (clk), .rst (rst), .g_input ({g_input[256], g_input[257], g_input[284], g_input[286], g_input[312]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[238]));
    dotproduct5 operation_conv239(.clk (clk), .rst (rst), .g_input ({g_input[257], g_input[258], g_input[285], g_input[287], g_input[313]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[239]));
    dotproduct5 operation_conv240(.clk (clk), .rst (rst), .g_input ({g_input[258], g_input[259], g_input[286], g_input[288], g_input[314]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[240]));
    dotproduct5 operation_conv241(.clk (clk), .rst (rst), .g_input ({g_input[259], g_input[260], g_input[287], g_input[289], g_input[315]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[241]));
    dotproduct5 operation_conv242(.clk (clk), .rst (rst), .g_input ({g_input[260], g_input[261], g_input[288], g_input[290], g_input[316]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[242]));
    dotproduct5 operation_conv243(.clk (clk), .rst (rst), .g_input ({g_input[261], g_input[262], g_input[289], g_input[291], g_input[317]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[243]));
    dotproduct5 operation_conv244(.clk (clk), .rst (rst), .g_input ({g_input[262], g_input[263], g_input[290], g_input[292], g_input[318]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[244]));
    dotproduct5 operation_conv245(.clk (clk), .rst (rst), .g_input ({g_input[263], g_input[264], g_input[291], g_input[293], g_input[319]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[245]));
    dotproduct5 operation_conv246(.clk (clk), .rst (rst), .g_input ({g_input[264], g_input[265], g_input[292], g_input[294], g_input[320]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[246]));
    dotproduct5 operation_conv247(.clk (clk), .rst (rst), .g_input ({g_input[265], g_input[266], g_input[293], g_input[295], g_input[321]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[247]));
    dotproduct5 operation_conv248(.clk (clk), .rst (rst), .g_input ({g_input[266], g_input[267], g_input[294], g_input[296], g_input[322]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[248]));
    dotproduct5 operation_conv249(.clk (clk), .rst (rst), .g_input ({g_input[267], g_input[268], g_input[295], g_input[297], g_input[323]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[249]));
    dotproduct5 operation_conv250(.clk (clk), .rst (rst), .g_input ({g_input[268], g_input[269], g_input[296], g_input[298], g_input[324]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[250]));
    dotproduct5 operation_conv251(.clk (clk), .rst (rst), .g_input ({g_input[269], g_input[270], g_input[297], g_input[299], g_input[325]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[251]));
    dotproduct5 operation_conv252(.clk (clk), .rst (rst), .g_input ({g_input[270], g_input[271], g_input[298], g_input[300], g_input[326]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[252]));
    dotproduct5 operation_conv253(.clk (clk), .rst (rst), .g_input ({g_input[271], g_input[272], g_input[299], g_input[301], g_input[327]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[253]));
    dotproduct5 operation_conv254(.clk (clk), .rst (rst), .g_input ({g_input[272], g_input[273], g_input[300], g_input[302], g_input[328]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[254]));
    dotproduct5 operation_conv255(.clk (clk), .rst (rst), .g_input ({g_input[273], g_input[274], g_input[301], g_input[303], g_input[329]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[255]));
    dotproduct5 operation_conv256(.clk (clk), .rst (rst), .g_input ({g_input[274], g_input[275], g_input[302], g_input[304], g_input[330]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[256]));
    dotproduct5 operation_conv257(.clk (clk), .rst (rst), .g_input ({g_input[275], g_input[276], g_input[303], g_input[305], g_input[331]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[257]));
    dotproduct5 operation_conv258(.clk (clk), .rst (rst), .g_input ({g_input[276], g_input[277], g_input[304], g_input[306], g_input[332]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[258]));
    dotproduct5 operation_conv259(.clk (clk), .rst (rst), .g_input ({g_input[277], g_input[278], g_input[305], g_input[307], g_input[333]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[259]));
    dotproduct5 operation_conv260(.clk (clk), .rst (rst), .g_input ({g_input[280], g_input[281], g_input[308], g_input[310], g_input[336]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[260]));
    dotproduct5 operation_conv261(.clk (clk), .rst (rst), .g_input ({g_input[281], g_input[282], g_input[309], g_input[311], g_input[337]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[261]));
    dotproduct5 operation_conv262(.clk (clk), .rst (rst), .g_input ({g_input[282], g_input[283], g_input[310], g_input[312], g_input[338]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[262]));
    dotproduct5 operation_conv263(.clk (clk), .rst (rst), .g_input ({g_input[283], g_input[284], g_input[311], g_input[313], g_input[339]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[263]));
    dotproduct5 operation_conv264(.clk (clk), .rst (rst), .g_input ({g_input[284], g_input[285], g_input[312], g_input[314], g_input[340]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[264]));
    dotproduct5 operation_conv265(.clk (clk), .rst (rst), .g_input ({g_input[285], g_input[286], g_input[313], g_input[315], g_input[341]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[265]));
    dotproduct5 operation_conv266(.clk (clk), .rst (rst), .g_input ({g_input[286], g_input[287], g_input[314], g_input[316], g_input[342]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[266]));
    dotproduct5 operation_conv267(.clk (clk), .rst (rst), .g_input ({g_input[287], g_input[288], g_input[315], g_input[317], g_input[343]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[267]));
    dotproduct5 operation_conv268(.clk (clk), .rst (rst), .g_input ({g_input[288], g_input[289], g_input[316], g_input[318], g_input[344]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[268]));
    dotproduct5 operation_conv269(.clk (clk), .rst (rst), .g_input ({g_input[289], g_input[290], g_input[317], g_input[319], g_input[345]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[269]));
    dotproduct5 operation_conv270(.clk (clk), .rst (rst), .g_input ({g_input[290], g_input[291], g_input[318], g_input[320], g_input[346]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[270]));
    dotproduct5 operation_conv271(.clk (clk), .rst (rst), .g_input ({g_input[291], g_input[292], g_input[319], g_input[321], g_input[347]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[271]));
    dotproduct5 operation_conv272(.clk (clk), .rst (rst), .g_input ({g_input[292], g_input[293], g_input[320], g_input[322], g_input[348]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[272]));
    dotproduct5 operation_conv273(.clk (clk), .rst (rst), .g_input ({g_input[293], g_input[294], g_input[321], g_input[323], g_input[349]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[273]));
    dotproduct5 operation_conv274(.clk (clk), .rst (rst), .g_input ({g_input[294], g_input[295], g_input[322], g_input[324], g_input[350]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[274]));
    dotproduct5 operation_conv275(.clk (clk), .rst (rst), .g_input ({g_input[295], g_input[296], g_input[323], g_input[325], g_input[351]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[275]));
    dotproduct5 operation_conv276(.clk (clk), .rst (rst), .g_input ({g_input[296], g_input[297], g_input[324], g_input[326], g_input[352]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[276]));
    dotproduct5 operation_conv277(.clk (clk), .rst (rst), .g_input ({g_input[297], g_input[298], g_input[325], g_input[327], g_input[353]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[277]));
    dotproduct5 operation_conv278(.clk (clk), .rst (rst), .g_input ({g_input[298], g_input[299], g_input[326], g_input[328], g_input[354]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[278]));
    dotproduct5 operation_conv279(.clk (clk), .rst (rst), .g_input ({g_input[299], g_input[300], g_input[327], g_input[329], g_input[355]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[279]));
    dotproduct5 operation_conv280(.clk (clk), .rst (rst), .g_input ({g_input[300], g_input[301], g_input[328], g_input[330], g_input[356]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[280]));
    dotproduct5 operation_conv281(.clk (clk), .rst (rst), .g_input ({g_input[301], g_input[302], g_input[329], g_input[331], g_input[357]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[281]));
    dotproduct5 operation_conv282(.clk (clk), .rst (rst), .g_input ({g_input[302], g_input[303], g_input[330], g_input[332], g_input[358]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[282]));
    dotproduct5 operation_conv283(.clk (clk), .rst (rst), .g_input ({g_input[303], g_input[304], g_input[331], g_input[333], g_input[359]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[283]));
    dotproduct5 operation_conv284(.clk (clk), .rst (rst), .g_input ({g_input[304], g_input[305], g_input[332], g_input[334], g_input[360]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[284]));
    dotproduct5 operation_conv285(.clk (clk), .rst (rst), .g_input ({g_input[305], g_input[306], g_input[333], g_input[335], g_input[361]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[285]));
    dotproduct5 operation_conv286(.clk (clk), .rst (rst), .g_input ({g_input[308], g_input[309], g_input[336], g_input[338], g_input[364]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[286]));
    dotproduct5 operation_conv287(.clk (clk), .rst (rst), .g_input ({g_input[309], g_input[310], g_input[337], g_input[339], g_input[365]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[287]));
    dotproduct5 operation_conv288(.clk (clk), .rst (rst), .g_input ({g_input[310], g_input[311], g_input[338], g_input[340], g_input[366]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[288]));
    dotproduct5 operation_conv289(.clk (clk), .rst (rst), .g_input ({g_input[311], g_input[312], g_input[339], g_input[341], g_input[367]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[289]));
    dotproduct5 operation_conv290(.clk (clk), .rst (rst), .g_input ({g_input[312], g_input[313], g_input[340], g_input[342], g_input[368]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[290]));
    dotproduct5 operation_conv291(.clk (clk), .rst (rst), .g_input ({g_input[313], g_input[314], g_input[341], g_input[343], g_input[369]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[291]));
    dotproduct5 operation_conv292(.clk (clk), .rst (rst), .g_input ({g_input[314], g_input[315], g_input[342], g_input[344], g_input[370]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[292]));
    dotproduct5 operation_conv293(.clk (clk), .rst (rst), .g_input ({g_input[315], g_input[316], g_input[343], g_input[345], g_input[371]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[293]));
    dotproduct5 operation_conv294(.clk (clk), .rst (rst), .g_input ({g_input[316], g_input[317], g_input[344], g_input[346], g_input[372]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[294]));
    dotproduct5 operation_conv295(.clk (clk), .rst (rst), .g_input ({g_input[317], g_input[318], g_input[345], g_input[347], g_input[373]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[295]));
    dotproduct5 operation_conv296(.clk (clk), .rst (rst), .g_input ({g_input[318], g_input[319], g_input[346], g_input[348], g_input[374]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[296]));
    dotproduct5 operation_conv297(.clk (clk), .rst (rst), .g_input ({g_input[319], g_input[320], g_input[347], g_input[349], g_input[375]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[297]));
    dotproduct5 operation_conv298(.clk (clk), .rst (rst), .g_input ({g_input[320], g_input[321], g_input[348], g_input[350], g_input[376]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[298]));
    dotproduct5 operation_conv299(.clk (clk), .rst (rst), .g_input ({g_input[321], g_input[322], g_input[349], g_input[351], g_input[377]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[299]));
    dotproduct5 operation_conv300(.clk (clk), .rst (rst), .g_input ({g_input[322], g_input[323], g_input[350], g_input[352], g_input[378]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[300]));
    dotproduct5 operation_conv301(.clk (clk), .rst (rst), .g_input ({g_input[323], g_input[324], g_input[351], g_input[353], g_input[379]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[301]));
    dotproduct5 operation_conv302(.clk (clk), .rst (rst), .g_input ({g_input[324], g_input[325], g_input[352], g_input[354], g_input[380]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[302]));
    dotproduct5 operation_conv303(.clk (clk), .rst (rst), .g_input ({g_input[325], g_input[326], g_input[353], g_input[355], g_input[381]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[303]));
    dotproduct5 operation_conv304(.clk (clk), .rst (rst), .g_input ({g_input[326], g_input[327], g_input[354], g_input[356], g_input[382]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[304]));
    dotproduct5 operation_conv305(.clk (clk), .rst (rst), .g_input ({g_input[327], g_input[328], g_input[355], g_input[357], g_input[383]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[305]));
    dotproduct5 operation_conv306(.clk (clk), .rst (rst), .g_input ({g_input[328], g_input[329], g_input[356], g_input[358], g_input[384]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[306]));
    dotproduct5 operation_conv307(.clk (clk), .rst (rst), .g_input ({g_input[329], g_input[330], g_input[357], g_input[359], g_input[385]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[307]));
    dotproduct5 operation_conv308(.clk (clk), .rst (rst), .g_input ({g_input[330], g_input[331], g_input[358], g_input[360], g_input[386]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[308]));
    dotproduct5 operation_conv309(.clk (clk), .rst (rst), .g_input ({g_input[331], g_input[332], g_input[359], g_input[361], g_input[387]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[309]));
    dotproduct5 operation_conv310(.clk (clk), .rst (rst), .g_input ({g_input[332], g_input[333], g_input[360], g_input[362], g_input[388]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[310]));
    dotproduct5 operation_conv311(.clk (clk), .rst (rst), .g_input ({g_input[333], g_input[334], g_input[361], g_input[363], g_input[389]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[311]));
    dotproduct5 operation_conv312(.clk (clk), .rst (rst), .g_input ({g_input[336], g_input[337], g_input[364], g_input[366], g_input[392]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[312]));
    dotproduct5 operation_conv313(.clk (clk), .rst (rst), .g_input ({g_input[337], g_input[338], g_input[365], g_input[367], g_input[393]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[313]));
    dotproduct5 operation_conv314(.clk (clk), .rst (rst), .g_input ({g_input[338], g_input[339], g_input[366], g_input[368], g_input[394]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[314]));
    dotproduct5 operation_conv315(.clk (clk), .rst (rst), .g_input ({g_input[339], g_input[340], g_input[367], g_input[369], g_input[395]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[315]));
    dotproduct5 operation_conv316(.clk (clk), .rst (rst), .g_input ({g_input[340], g_input[341], g_input[368], g_input[370], g_input[396]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[316]));
    dotproduct5 operation_conv317(.clk (clk), .rst (rst), .g_input ({g_input[341], g_input[342], g_input[369], g_input[371], g_input[397]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[317]));
    dotproduct5 operation_conv318(.clk (clk), .rst (rst), .g_input ({g_input[342], g_input[343], g_input[370], g_input[372], g_input[398]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[318]));
    dotproduct5 operation_conv319(.clk (clk), .rst (rst), .g_input ({g_input[343], g_input[344], g_input[371], g_input[373], g_input[399]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[319]));
    dotproduct5 operation_conv320(.clk (clk), .rst (rst), .g_input ({g_input[344], g_input[345], g_input[372], g_input[374], g_input[400]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[320]));
    dotproduct5 operation_conv321(.clk (clk), .rst (rst), .g_input ({g_input[345], g_input[346], g_input[373], g_input[375], g_input[401]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[321]));
    dotproduct5 operation_conv322(.clk (clk), .rst (rst), .g_input ({g_input[346], g_input[347], g_input[374], g_input[376], g_input[402]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[322]));
    dotproduct5 operation_conv323(.clk (clk), .rst (rst), .g_input ({g_input[347], g_input[348], g_input[375], g_input[377], g_input[403]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[323]));
    dotproduct5 operation_conv324(.clk (clk), .rst (rst), .g_input ({g_input[348], g_input[349], g_input[376], g_input[378], g_input[404]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[324]));
    dotproduct5 operation_conv325(.clk (clk), .rst (rst), .g_input ({g_input[349], g_input[350], g_input[377], g_input[379], g_input[405]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[325]));
    dotproduct5 operation_conv326(.clk (clk), .rst (rst), .g_input ({g_input[350], g_input[351], g_input[378], g_input[380], g_input[406]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[326]));
    dotproduct5 operation_conv327(.clk (clk), .rst (rst), .g_input ({g_input[351], g_input[352], g_input[379], g_input[381], g_input[407]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[327]));
    dotproduct5 operation_conv328(.clk (clk), .rst (rst), .g_input ({g_input[352], g_input[353], g_input[380], g_input[382], g_input[408]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[328]));
    dotproduct5 operation_conv329(.clk (clk), .rst (rst), .g_input ({g_input[353], g_input[354], g_input[381], g_input[383], g_input[409]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[329]));
    dotproduct5 operation_conv330(.clk (clk), .rst (rst), .g_input ({g_input[354], g_input[355], g_input[382], g_input[384], g_input[410]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[330]));
    dotproduct5 operation_conv331(.clk (clk), .rst (rst), .g_input ({g_input[355], g_input[356], g_input[383], g_input[385], g_input[411]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[331]));
    dotproduct5 operation_conv332(.clk (clk), .rst (rst), .g_input ({g_input[356], g_input[357], g_input[384], g_input[386], g_input[412]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[332]));
    dotproduct5 operation_conv333(.clk (clk), .rst (rst), .g_input ({g_input[357], g_input[358], g_input[385], g_input[387], g_input[413]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[333]));
    dotproduct5 operation_conv334(.clk (clk), .rst (rst), .g_input ({g_input[358], g_input[359], g_input[386], g_input[388], g_input[414]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[334]));
    dotproduct5 operation_conv335(.clk (clk), .rst (rst), .g_input ({g_input[359], g_input[360], g_input[387], g_input[389], g_input[415]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[335]));
    dotproduct5 operation_conv336(.clk (clk), .rst (rst), .g_input ({g_input[360], g_input[361], g_input[388], g_input[390], g_input[416]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[336]));
    dotproduct5 operation_conv337(.clk (clk), .rst (rst), .g_input ({g_input[361], g_input[362], g_input[389], g_input[391], g_input[417]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[337]));
    dotproduct5 operation_conv338(.clk (clk), .rst (rst), .g_input ({g_input[364], g_input[365], g_input[392], g_input[394], g_input[420]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[338]));
    dotproduct5 operation_conv339(.clk (clk), .rst (rst), .g_input ({g_input[365], g_input[366], g_input[393], g_input[395], g_input[421]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[339]));
    dotproduct5 operation_conv340(.clk (clk), .rst (rst), .g_input ({g_input[366], g_input[367], g_input[394], g_input[396], g_input[422]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[340]));
    dotproduct5 operation_conv341(.clk (clk), .rst (rst), .g_input ({g_input[367], g_input[368], g_input[395], g_input[397], g_input[423]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[341]));
    dotproduct5 operation_conv342(.clk (clk), .rst (rst), .g_input ({g_input[368], g_input[369], g_input[396], g_input[398], g_input[424]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[342]));
    dotproduct5 operation_conv343(.clk (clk), .rst (rst), .g_input ({g_input[369], g_input[370], g_input[397], g_input[399], g_input[425]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[343]));
    dotproduct5 operation_conv344(.clk (clk), .rst (rst), .g_input ({g_input[370], g_input[371], g_input[398], g_input[400], g_input[426]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[344]));
    dotproduct5 operation_conv345(.clk (clk), .rst (rst), .g_input ({g_input[371], g_input[372], g_input[399], g_input[401], g_input[427]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[345]));
    dotproduct5 operation_conv346(.clk (clk), .rst (rst), .g_input ({g_input[372], g_input[373], g_input[400], g_input[402], g_input[428]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[346]));
    dotproduct5 operation_conv347(.clk (clk), .rst (rst), .g_input ({g_input[373], g_input[374], g_input[401], g_input[403], g_input[429]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[347]));
    dotproduct5 operation_conv348(.clk (clk), .rst (rst), .g_input ({g_input[374], g_input[375], g_input[402], g_input[404], g_input[430]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[348]));
    dotproduct5 operation_conv349(.clk (clk), .rst (rst), .g_input ({g_input[375], g_input[376], g_input[403], g_input[405], g_input[431]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[349]));
    dotproduct5 operation_conv350(.clk (clk), .rst (rst), .g_input ({g_input[376], g_input[377], g_input[404], g_input[406], g_input[432]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[350]));
    dotproduct5 operation_conv351(.clk (clk), .rst (rst), .g_input ({g_input[377], g_input[378], g_input[405], g_input[407], g_input[433]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[351]));
    dotproduct5 operation_conv352(.clk (clk), .rst (rst), .g_input ({g_input[378], g_input[379], g_input[406], g_input[408], g_input[434]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[352]));
    dotproduct5 operation_conv353(.clk (clk), .rst (rst), .g_input ({g_input[379], g_input[380], g_input[407], g_input[409], g_input[435]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[353]));
    dotproduct5 operation_conv354(.clk (clk), .rst (rst), .g_input ({g_input[380], g_input[381], g_input[408], g_input[410], g_input[436]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[354]));
    dotproduct5 operation_conv355(.clk (clk), .rst (rst), .g_input ({g_input[381], g_input[382], g_input[409], g_input[411], g_input[437]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[355]));
    dotproduct5 operation_conv356(.clk (clk), .rst (rst), .g_input ({g_input[382], g_input[383], g_input[410], g_input[412], g_input[438]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[356]));
    dotproduct5 operation_conv357(.clk (clk), .rst (rst), .g_input ({g_input[383], g_input[384], g_input[411], g_input[413], g_input[439]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[357]));
    dotproduct5 operation_conv358(.clk (clk), .rst (rst), .g_input ({g_input[384], g_input[385], g_input[412], g_input[414], g_input[440]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[358]));
    dotproduct5 operation_conv359(.clk (clk), .rst (rst), .g_input ({g_input[385], g_input[386], g_input[413], g_input[415], g_input[441]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[359]));
    dotproduct5 operation_conv360(.clk (clk), .rst (rst), .g_input ({g_input[386], g_input[387], g_input[414], g_input[416], g_input[442]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[360]));
    dotproduct5 operation_conv361(.clk (clk), .rst (rst), .g_input ({g_input[387], g_input[388], g_input[415], g_input[417], g_input[443]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[361]));
    dotproduct5 operation_conv362(.clk (clk), .rst (rst), .g_input ({g_input[388], g_input[389], g_input[416], g_input[418], g_input[444]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[362]));
    dotproduct5 operation_conv363(.clk (clk), .rst (rst), .g_input ({g_input[389], g_input[390], g_input[417], g_input[419], g_input[445]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[363]));
    dotproduct5 operation_conv364(.clk (clk), .rst (rst), .g_input ({g_input[392], g_input[393], g_input[420], g_input[422], g_input[448]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[364]));
    dotproduct5 operation_conv365(.clk (clk), .rst (rst), .g_input ({g_input[393], g_input[394], g_input[421], g_input[423], g_input[449]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[365]));
    dotproduct5 operation_conv366(.clk (clk), .rst (rst), .g_input ({g_input[394], g_input[395], g_input[422], g_input[424], g_input[450]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[366]));
    dotproduct5 operation_conv367(.clk (clk), .rst (rst), .g_input ({g_input[395], g_input[396], g_input[423], g_input[425], g_input[451]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[367]));
    dotproduct5 operation_conv368(.clk (clk), .rst (rst), .g_input ({g_input[396], g_input[397], g_input[424], g_input[426], g_input[452]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[368]));
    dotproduct5 operation_conv369(.clk (clk), .rst (rst), .g_input ({g_input[397], g_input[398], g_input[425], g_input[427], g_input[453]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[369]));
    dotproduct5 operation_conv370(.clk (clk), .rst (rst), .g_input ({g_input[398], g_input[399], g_input[426], g_input[428], g_input[454]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[370]));
    dotproduct5 operation_conv371(.clk (clk), .rst (rst), .g_input ({g_input[399], g_input[400], g_input[427], g_input[429], g_input[455]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[371]));
    dotproduct5 operation_conv372(.clk (clk), .rst (rst), .g_input ({g_input[400], g_input[401], g_input[428], g_input[430], g_input[456]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[372]));
    dotproduct5 operation_conv373(.clk (clk), .rst (rst), .g_input ({g_input[401], g_input[402], g_input[429], g_input[431], g_input[457]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[373]));
    dotproduct5 operation_conv374(.clk (clk), .rst (rst), .g_input ({g_input[402], g_input[403], g_input[430], g_input[432], g_input[458]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[374]));
    dotproduct5 operation_conv375(.clk (clk), .rst (rst), .g_input ({g_input[403], g_input[404], g_input[431], g_input[433], g_input[459]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[375]));
    dotproduct5 operation_conv376(.clk (clk), .rst (rst), .g_input ({g_input[404], g_input[405], g_input[432], g_input[434], g_input[460]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[376]));
    dotproduct5 operation_conv377(.clk (clk), .rst (rst), .g_input ({g_input[405], g_input[406], g_input[433], g_input[435], g_input[461]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[377]));
    dotproduct5 operation_conv378(.clk (clk), .rst (rst), .g_input ({g_input[406], g_input[407], g_input[434], g_input[436], g_input[462]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[378]));
    dotproduct5 operation_conv379(.clk (clk), .rst (rst), .g_input ({g_input[407], g_input[408], g_input[435], g_input[437], g_input[463]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[379]));
    dotproduct5 operation_conv380(.clk (clk), .rst (rst), .g_input ({g_input[408], g_input[409], g_input[436], g_input[438], g_input[464]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[380]));
    dotproduct5 operation_conv381(.clk (clk), .rst (rst), .g_input ({g_input[409], g_input[410], g_input[437], g_input[439], g_input[465]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[381]));
    dotproduct5 operation_conv382(.clk (clk), .rst (rst), .g_input ({g_input[410], g_input[411], g_input[438], g_input[440], g_input[466]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[382]));
    dotproduct5 operation_conv383(.clk (clk), .rst (rst), .g_input ({g_input[411], g_input[412], g_input[439], g_input[441], g_input[467]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[383]));
    dotproduct5 operation_conv384(.clk (clk), .rst (rst), .g_input ({g_input[412], g_input[413], g_input[440], g_input[442], g_input[468]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[384]));
    dotproduct5 operation_conv385(.clk (clk), .rst (rst), .g_input ({g_input[413], g_input[414], g_input[441], g_input[443], g_input[469]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[385]));
    dotproduct5 operation_conv386(.clk (clk), .rst (rst), .g_input ({g_input[414], g_input[415], g_input[442], g_input[444], g_input[470]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[386]));
    dotproduct5 operation_conv387(.clk (clk), .rst (rst), .g_input ({g_input[415], g_input[416], g_input[443], g_input[445], g_input[471]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[387]));
    dotproduct5 operation_conv388(.clk (clk), .rst (rst), .g_input ({g_input[416], g_input[417], g_input[444], g_input[446], g_input[472]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[388]));
    dotproduct5 operation_conv389(.clk (clk), .rst (rst), .g_input ({g_input[417], g_input[418], g_input[445], g_input[447], g_input[473]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[389]));
    dotproduct5 operation_conv390(.clk (clk), .rst (rst), .g_input ({g_input[420], g_input[421], g_input[448], g_input[450], g_input[476]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[390]));
    dotproduct5 operation_conv391(.clk (clk), .rst (rst), .g_input ({g_input[421], g_input[422], g_input[449], g_input[451], g_input[477]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[391]));
    dotproduct5 operation_conv392(.clk (clk), .rst (rst), .g_input ({g_input[422], g_input[423], g_input[450], g_input[452], g_input[478]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[392]));
    dotproduct5 operation_conv393(.clk (clk), .rst (rst), .g_input ({g_input[423], g_input[424], g_input[451], g_input[453], g_input[479]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[393]));
    dotproduct5 operation_conv394(.clk (clk), .rst (rst), .g_input ({g_input[424], g_input[425], g_input[452], g_input[454], g_input[480]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[394]));
    dotproduct5 operation_conv395(.clk (clk), .rst (rst), .g_input ({g_input[425], g_input[426], g_input[453], g_input[455], g_input[481]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[395]));
    dotproduct5 operation_conv396(.clk (clk), .rst (rst), .g_input ({g_input[426], g_input[427], g_input[454], g_input[456], g_input[482]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[396]));
    dotproduct5 operation_conv397(.clk (clk), .rst (rst), .g_input ({g_input[427], g_input[428], g_input[455], g_input[457], g_input[483]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[397]));
    dotproduct5 operation_conv398(.clk (clk), .rst (rst), .g_input ({g_input[428], g_input[429], g_input[456], g_input[458], g_input[484]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[398]));
    dotproduct5 operation_conv399(.clk (clk), .rst (rst), .g_input ({g_input[429], g_input[430], g_input[457], g_input[459], g_input[485]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[399]));
    dotproduct5 operation_conv400(.clk (clk), .rst (rst), .g_input ({g_input[430], g_input[431], g_input[458], g_input[460], g_input[486]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[400]));
    dotproduct5 operation_conv401(.clk (clk), .rst (rst), .g_input ({g_input[431], g_input[432], g_input[459], g_input[461], g_input[487]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[401]));
    dotproduct5 operation_conv402(.clk (clk), .rst (rst), .g_input ({g_input[432], g_input[433], g_input[460], g_input[462], g_input[488]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[402]));
    dotproduct5 operation_conv403(.clk (clk), .rst (rst), .g_input ({g_input[433], g_input[434], g_input[461], g_input[463], g_input[489]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[403]));
    dotproduct5 operation_conv404(.clk (clk), .rst (rst), .g_input ({g_input[434], g_input[435], g_input[462], g_input[464], g_input[490]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[404]));
    dotproduct5 operation_conv405(.clk (clk), .rst (rst), .g_input ({g_input[435], g_input[436], g_input[463], g_input[465], g_input[491]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[405]));
    dotproduct5 operation_conv406(.clk (clk), .rst (rst), .g_input ({g_input[436], g_input[437], g_input[464], g_input[466], g_input[492]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[406]));
    dotproduct5 operation_conv407(.clk (clk), .rst (rst), .g_input ({g_input[437], g_input[438], g_input[465], g_input[467], g_input[493]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[407]));
    dotproduct5 operation_conv408(.clk (clk), .rst (rst), .g_input ({g_input[438], g_input[439], g_input[466], g_input[468], g_input[494]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[408]));
    dotproduct5 operation_conv409(.clk (clk), .rst (rst), .g_input ({g_input[439], g_input[440], g_input[467], g_input[469], g_input[495]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[409]));
    dotproduct5 operation_conv410(.clk (clk), .rst (rst), .g_input ({g_input[440], g_input[441], g_input[468], g_input[470], g_input[496]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[410]));
    dotproduct5 operation_conv411(.clk (clk), .rst (rst), .g_input ({g_input[441], g_input[442], g_input[469], g_input[471], g_input[497]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[411]));
    dotproduct5 operation_conv412(.clk (clk), .rst (rst), .g_input ({g_input[442], g_input[443], g_input[470], g_input[472], g_input[498]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[412]));
    dotproduct5 operation_conv413(.clk (clk), .rst (rst), .g_input ({g_input[443], g_input[444], g_input[471], g_input[473], g_input[499]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[413]));
    dotproduct5 operation_conv414(.clk (clk), .rst (rst), .g_input ({g_input[444], g_input[445], g_input[472], g_input[474], g_input[500]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[414]));
    dotproduct5 operation_conv415(.clk (clk), .rst (rst), .g_input ({g_input[445], g_input[446], g_input[473], g_input[475], g_input[501]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[415]));
    dotproduct5 operation_conv416(.clk (clk), .rst (rst), .g_input ({g_input[448], g_input[449], g_input[476], g_input[478], g_input[504]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[416]));
    dotproduct5 operation_conv417(.clk (clk), .rst (rst), .g_input ({g_input[449], g_input[450], g_input[477], g_input[479], g_input[505]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[417]));
    dotproduct5 operation_conv418(.clk (clk), .rst (rst), .g_input ({g_input[450], g_input[451], g_input[478], g_input[480], g_input[506]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[418]));
    dotproduct5 operation_conv419(.clk (clk), .rst (rst), .g_input ({g_input[451], g_input[452], g_input[479], g_input[481], g_input[507]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[419]));
    dotproduct5 operation_conv420(.clk (clk), .rst (rst), .g_input ({g_input[452], g_input[453], g_input[480], g_input[482], g_input[508]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[420]));
    dotproduct5 operation_conv421(.clk (clk), .rst (rst), .g_input ({g_input[453], g_input[454], g_input[481], g_input[483], g_input[509]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[421]));
    dotproduct5 operation_conv422(.clk (clk), .rst (rst), .g_input ({g_input[454], g_input[455], g_input[482], g_input[484], g_input[510]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[422]));
    dotproduct5 operation_conv423(.clk (clk), .rst (rst), .g_input ({g_input[455], g_input[456], g_input[483], g_input[485], g_input[511]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[423]));
    dotproduct5 operation_conv424(.clk (clk), .rst (rst), .g_input ({g_input[456], g_input[457], g_input[484], g_input[486], g_input[512]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[424]));
    dotproduct5 operation_conv425(.clk (clk), .rst (rst), .g_input ({g_input[457], g_input[458], g_input[485], g_input[487], g_input[513]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[425]));
    dotproduct5 operation_conv426(.clk (clk), .rst (rst), .g_input ({g_input[458], g_input[459], g_input[486], g_input[488], g_input[514]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[426]));
    dotproduct5 operation_conv427(.clk (clk), .rst (rst), .g_input ({g_input[459], g_input[460], g_input[487], g_input[489], g_input[515]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[427]));
    dotproduct5 operation_conv428(.clk (clk), .rst (rst), .g_input ({g_input[460], g_input[461], g_input[488], g_input[490], g_input[516]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[428]));
    dotproduct5 operation_conv429(.clk (clk), .rst (rst), .g_input ({g_input[461], g_input[462], g_input[489], g_input[491], g_input[517]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[429]));
    dotproduct5 operation_conv430(.clk (clk), .rst (rst), .g_input ({g_input[462], g_input[463], g_input[490], g_input[492], g_input[518]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[430]));
    dotproduct5 operation_conv431(.clk (clk), .rst (rst), .g_input ({g_input[463], g_input[464], g_input[491], g_input[493], g_input[519]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[431]));
    dotproduct5 operation_conv432(.clk (clk), .rst (rst), .g_input ({g_input[464], g_input[465], g_input[492], g_input[494], g_input[520]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[432]));
    dotproduct5 operation_conv433(.clk (clk), .rst (rst), .g_input ({g_input[465], g_input[466], g_input[493], g_input[495], g_input[521]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[433]));
    dotproduct5 operation_conv434(.clk (clk), .rst (rst), .g_input ({g_input[466], g_input[467], g_input[494], g_input[496], g_input[522]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[434]));
    dotproduct5 operation_conv435(.clk (clk), .rst (rst), .g_input ({g_input[467], g_input[468], g_input[495], g_input[497], g_input[523]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[435]));
    dotproduct5 operation_conv436(.clk (clk), .rst (rst), .g_input ({g_input[468], g_input[469], g_input[496], g_input[498], g_input[524]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[436]));
    dotproduct5 operation_conv437(.clk (clk), .rst (rst), .g_input ({g_input[469], g_input[470], g_input[497], g_input[499], g_input[525]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[437]));
    dotproduct5 operation_conv438(.clk (clk), .rst (rst), .g_input ({g_input[470], g_input[471], g_input[498], g_input[500], g_input[526]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[438]));
    dotproduct5 operation_conv439(.clk (clk), .rst (rst), .g_input ({g_input[471], g_input[472], g_input[499], g_input[501], g_input[527]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[439]));
    dotproduct5 operation_conv440(.clk (clk), .rst (rst), .g_input ({g_input[472], g_input[473], g_input[500], g_input[502], g_input[528]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[440]));
    dotproduct5 operation_conv441(.clk (clk), .rst (rst), .g_input ({g_input[473], g_input[474], g_input[501], g_input[503], g_input[529]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[441]));
    dotproduct5 operation_conv442(.clk (clk), .rst (rst), .g_input ({g_input[476], g_input[477], g_input[504], g_input[506], g_input[532]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[442]));
    dotproduct5 operation_conv443(.clk (clk), .rst (rst), .g_input ({g_input[477], g_input[478], g_input[505], g_input[507], g_input[533]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[443]));
    dotproduct5 operation_conv444(.clk (clk), .rst (rst), .g_input ({g_input[478], g_input[479], g_input[506], g_input[508], g_input[534]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[444]));
    dotproduct5 operation_conv445(.clk (clk), .rst (rst), .g_input ({g_input[479], g_input[480], g_input[507], g_input[509], g_input[535]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[445]));
    dotproduct5 operation_conv446(.clk (clk), .rst (rst), .g_input ({g_input[480], g_input[481], g_input[508], g_input[510], g_input[536]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[446]));
    dotproduct5 operation_conv447(.clk (clk), .rst (rst), .g_input ({g_input[481], g_input[482], g_input[509], g_input[511], g_input[537]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[447]));
    dotproduct5 operation_conv448(.clk (clk), .rst (rst), .g_input ({g_input[482], g_input[483], g_input[510], g_input[512], g_input[538]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[448]));
    dotproduct5 operation_conv449(.clk (clk), .rst (rst), .g_input ({g_input[483], g_input[484], g_input[511], g_input[513], g_input[539]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[449]));
    dotproduct5 operation_conv450(.clk (clk), .rst (rst), .g_input ({g_input[484], g_input[485], g_input[512], g_input[514], g_input[540]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[450]));
    dotproduct5 operation_conv451(.clk (clk), .rst (rst), .g_input ({g_input[485], g_input[486], g_input[513], g_input[515], g_input[541]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[451]));
    dotproduct5 operation_conv452(.clk (clk), .rst (rst), .g_input ({g_input[486], g_input[487], g_input[514], g_input[516], g_input[542]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[452]));
    dotproduct5 operation_conv453(.clk (clk), .rst (rst), .g_input ({g_input[487], g_input[488], g_input[515], g_input[517], g_input[543]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[453]));
    dotproduct5 operation_conv454(.clk (clk), .rst (rst), .g_input ({g_input[488], g_input[489], g_input[516], g_input[518], g_input[544]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[454]));
    dotproduct5 operation_conv455(.clk (clk), .rst (rst), .g_input ({g_input[489], g_input[490], g_input[517], g_input[519], g_input[545]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[455]));
    dotproduct5 operation_conv456(.clk (clk), .rst (rst), .g_input ({g_input[490], g_input[491], g_input[518], g_input[520], g_input[546]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[456]));
    dotproduct5 operation_conv457(.clk (clk), .rst (rst), .g_input ({g_input[491], g_input[492], g_input[519], g_input[521], g_input[547]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[457]));
    dotproduct5 operation_conv458(.clk (clk), .rst (rst), .g_input ({g_input[492], g_input[493], g_input[520], g_input[522], g_input[548]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[458]));
    dotproduct5 operation_conv459(.clk (clk), .rst (rst), .g_input ({g_input[493], g_input[494], g_input[521], g_input[523], g_input[549]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[459]));
    dotproduct5 operation_conv460(.clk (clk), .rst (rst), .g_input ({g_input[494], g_input[495], g_input[522], g_input[524], g_input[550]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[460]));
    dotproduct5 operation_conv461(.clk (clk), .rst (rst), .g_input ({g_input[495], g_input[496], g_input[523], g_input[525], g_input[551]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[461]));
    dotproduct5 operation_conv462(.clk (clk), .rst (rst), .g_input ({g_input[496], g_input[497], g_input[524], g_input[526], g_input[552]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[462]));
    dotproduct5 operation_conv463(.clk (clk), .rst (rst), .g_input ({g_input[497], g_input[498], g_input[525], g_input[527], g_input[553]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[463]));
    dotproduct5 operation_conv464(.clk (clk), .rst (rst), .g_input ({g_input[498], g_input[499], g_input[526], g_input[528], g_input[554]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[464]));
    dotproduct5 operation_conv465(.clk (clk), .rst (rst), .g_input ({g_input[499], g_input[500], g_input[527], g_input[529], g_input[555]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[465]));
    dotproduct5 operation_conv466(.clk (clk), .rst (rst), .g_input ({g_input[500], g_input[501], g_input[528], g_input[530], g_input[556]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[466]));
    dotproduct5 operation_conv467(.clk (clk), .rst (rst), .g_input ({g_input[501], g_input[502], g_input[529], g_input[531], g_input[557]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[467]));
    dotproduct5 operation_conv468(.clk (clk), .rst (rst), .g_input ({g_input[504], g_input[505], g_input[532], g_input[534], g_input[560]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[468]));
    dotproduct5 operation_conv469(.clk (clk), .rst (rst), .g_input ({g_input[505], g_input[506], g_input[533], g_input[535], g_input[561]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[469]));
    dotproduct5 operation_conv470(.clk (clk), .rst (rst), .g_input ({g_input[506], g_input[507], g_input[534], g_input[536], g_input[562]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[470]));
    dotproduct5 operation_conv471(.clk (clk), .rst (rst), .g_input ({g_input[507], g_input[508], g_input[535], g_input[537], g_input[563]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[471]));
    dotproduct5 operation_conv472(.clk (clk), .rst (rst), .g_input ({g_input[508], g_input[509], g_input[536], g_input[538], g_input[564]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[472]));
    dotproduct5 operation_conv473(.clk (clk), .rst (rst), .g_input ({g_input[509], g_input[510], g_input[537], g_input[539], g_input[565]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[473]));
    dotproduct5 operation_conv474(.clk (clk), .rst (rst), .g_input ({g_input[510], g_input[511], g_input[538], g_input[540], g_input[566]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[474]));
    dotproduct5 operation_conv475(.clk (clk), .rst (rst), .g_input ({g_input[511], g_input[512], g_input[539], g_input[541], g_input[567]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[475]));
    dotproduct5 operation_conv476(.clk (clk), .rst (rst), .g_input ({g_input[512], g_input[513], g_input[540], g_input[542], g_input[568]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[476]));
    dotproduct5 operation_conv477(.clk (clk), .rst (rst), .g_input ({g_input[513], g_input[514], g_input[541], g_input[543], g_input[569]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[477]));
    dotproduct5 operation_conv478(.clk (clk), .rst (rst), .g_input ({g_input[514], g_input[515], g_input[542], g_input[544], g_input[570]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[478]));
    dotproduct5 operation_conv479(.clk (clk), .rst (rst), .g_input ({g_input[515], g_input[516], g_input[543], g_input[545], g_input[571]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[479]));
    dotproduct5 operation_conv480(.clk (clk), .rst (rst), .g_input ({g_input[516], g_input[517], g_input[544], g_input[546], g_input[572]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[480]));
    dotproduct5 operation_conv481(.clk (clk), .rst (rst), .g_input ({g_input[517], g_input[518], g_input[545], g_input[547], g_input[573]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[481]));
    dotproduct5 operation_conv482(.clk (clk), .rst (rst), .g_input ({g_input[518], g_input[519], g_input[546], g_input[548], g_input[574]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[482]));
    dotproduct5 operation_conv483(.clk (clk), .rst (rst), .g_input ({g_input[519], g_input[520], g_input[547], g_input[549], g_input[575]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[483]));
    dotproduct5 operation_conv484(.clk (clk), .rst (rst), .g_input ({g_input[520], g_input[521], g_input[548], g_input[550], g_input[576]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[484]));
    dotproduct5 operation_conv485(.clk (clk), .rst (rst), .g_input ({g_input[521], g_input[522], g_input[549], g_input[551], g_input[577]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[485]));
    dotproduct5 operation_conv486(.clk (clk), .rst (rst), .g_input ({g_input[522], g_input[523], g_input[550], g_input[552], g_input[578]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[486]));
    dotproduct5 operation_conv487(.clk (clk), .rst (rst), .g_input ({g_input[523], g_input[524], g_input[551], g_input[553], g_input[579]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[487]));
    dotproduct5 operation_conv488(.clk (clk), .rst (rst), .g_input ({g_input[524], g_input[525], g_input[552], g_input[554], g_input[580]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[488]));
    dotproduct5 operation_conv489(.clk (clk), .rst (rst), .g_input ({g_input[525], g_input[526], g_input[553], g_input[555], g_input[581]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[489]));
    dotproduct5 operation_conv490(.clk (clk), .rst (rst), .g_input ({g_input[526], g_input[527], g_input[554], g_input[556], g_input[582]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[490]));
    dotproduct5 operation_conv491(.clk (clk), .rst (rst), .g_input ({g_input[527], g_input[528], g_input[555], g_input[557], g_input[583]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[491]));
    dotproduct5 operation_conv492(.clk (clk), .rst (rst), .g_input ({g_input[528], g_input[529], g_input[556], g_input[558], g_input[584]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[492]));
    dotproduct5 operation_conv493(.clk (clk), .rst (rst), .g_input ({g_input[529], g_input[530], g_input[557], g_input[559], g_input[585]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[493]));
    dotproduct5 operation_conv494(.clk (clk), .rst (rst), .g_input ({g_input[532], g_input[533], g_input[560], g_input[562], g_input[588]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[494]));
    dotproduct5 operation_conv495(.clk (clk), .rst (rst), .g_input ({g_input[533], g_input[534], g_input[561], g_input[563], g_input[589]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[495]));
    dotproduct5 operation_conv496(.clk (clk), .rst (rst), .g_input ({g_input[534], g_input[535], g_input[562], g_input[564], g_input[590]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[496]));
    dotproduct5 operation_conv497(.clk (clk), .rst (rst), .g_input ({g_input[535], g_input[536], g_input[563], g_input[565], g_input[591]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[497]));
    dotproduct5 operation_conv498(.clk (clk), .rst (rst), .g_input ({g_input[536], g_input[537], g_input[564], g_input[566], g_input[592]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[498]));
    dotproduct5 operation_conv499(.clk (clk), .rst (rst), .g_input ({g_input[537], g_input[538], g_input[565], g_input[567], g_input[593]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[499]));
    dotproduct5 operation_conv500(.clk (clk), .rst (rst), .g_input ({g_input[538], g_input[539], g_input[566], g_input[568], g_input[594]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[500]));
    dotproduct5 operation_conv501(.clk (clk), .rst (rst), .g_input ({g_input[539], g_input[540], g_input[567], g_input[569], g_input[595]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[501]));
    dotproduct5 operation_conv502(.clk (clk), .rst (rst), .g_input ({g_input[540], g_input[541], g_input[568], g_input[570], g_input[596]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[502]));
    dotproduct5 operation_conv503(.clk (clk), .rst (rst), .g_input ({g_input[541], g_input[542], g_input[569], g_input[571], g_input[597]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[503]));
    dotproduct5 operation_conv504(.clk (clk), .rst (rst), .g_input ({g_input[542], g_input[543], g_input[570], g_input[572], g_input[598]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[504]));
    dotproduct5 operation_conv505(.clk (clk), .rst (rst), .g_input ({g_input[543], g_input[544], g_input[571], g_input[573], g_input[599]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[505]));
    dotproduct5 operation_conv506(.clk (clk), .rst (rst), .g_input ({g_input[544], g_input[545], g_input[572], g_input[574], g_input[600]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[506]));
    dotproduct5 operation_conv507(.clk (clk), .rst (rst), .g_input ({g_input[545], g_input[546], g_input[573], g_input[575], g_input[601]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[507]));
    dotproduct5 operation_conv508(.clk (clk), .rst (rst), .g_input ({g_input[546], g_input[547], g_input[574], g_input[576], g_input[602]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[508]));
    dotproduct5 operation_conv509(.clk (clk), .rst (rst), .g_input ({g_input[547], g_input[548], g_input[575], g_input[577], g_input[603]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[509]));
    dotproduct5 operation_conv510(.clk (clk), .rst (rst), .g_input ({g_input[548], g_input[549], g_input[576], g_input[578], g_input[604]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[510]));
    dotproduct5 operation_conv511(.clk (clk), .rst (rst), .g_input ({g_input[549], g_input[550], g_input[577], g_input[579], g_input[605]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[511]));
    dotproduct5 operation_conv512(.clk (clk), .rst (rst), .g_input ({g_input[550], g_input[551], g_input[578], g_input[580], g_input[606]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[512]));
    dotproduct5 operation_conv513(.clk (clk), .rst (rst), .g_input ({g_input[551], g_input[552], g_input[579], g_input[581], g_input[607]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[513]));
    dotproduct5 operation_conv514(.clk (clk), .rst (rst), .g_input ({g_input[552], g_input[553], g_input[580], g_input[582], g_input[608]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[514]));
    dotproduct5 operation_conv515(.clk (clk), .rst (rst), .g_input ({g_input[553], g_input[554], g_input[581], g_input[583], g_input[609]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[515]));
    dotproduct5 operation_conv516(.clk (clk), .rst (rst), .g_input ({g_input[554], g_input[555], g_input[582], g_input[584], g_input[610]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[516]));
    dotproduct5 operation_conv517(.clk (clk), .rst (rst), .g_input ({g_input[555], g_input[556], g_input[583], g_input[585], g_input[611]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[517]));
    dotproduct5 operation_conv518(.clk (clk), .rst (rst), .g_input ({g_input[556], g_input[557], g_input[584], g_input[586], g_input[612]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[518]));
    dotproduct5 operation_conv519(.clk (clk), .rst (rst), .g_input ({g_input[557], g_input[558], g_input[585], g_input[587], g_input[613]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[519]));
    dotproduct5 operation_conv520(.clk (clk), .rst (rst), .g_input ({g_input[560], g_input[561], g_input[588], g_input[590], g_input[616]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[520]));
    dotproduct5 operation_conv521(.clk (clk), .rst (rst), .g_input ({g_input[561], g_input[562], g_input[589], g_input[591], g_input[617]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[521]));
    dotproduct5 operation_conv522(.clk (clk), .rst (rst), .g_input ({g_input[562], g_input[563], g_input[590], g_input[592], g_input[618]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[522]));
    dotproduct5 operation_conv523(.clk (clk), .rst (rst), .g_input ({g_input[563], g_input[564], g_input[591], g_input[593], g_input[619]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[523]));
    dotproduct5 operation_conv524(.clk (clk), .rst (rst), .g_input ({g_input[564], g_input[565], g_input[592], g_input[594], g_input[620]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[524]));
    dotproduct5 operation_conv525(.clk (clk), .rst (rst), .g_input ({g_input[565], g_input[566], g_input[593], g_input[595], g_input[621]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[525]));
    dotproduct5 operation_conv526(.clk (clk), .rst (rst), .g_input ({g_input[566], g_input[567], g_input[594], g_input[596], g_input[622]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[526]));
    dotproduct5 operation_conv527(.clk (clk), .rst (rst), .g_input ({g_input[567], g_input[568], g_input[595], g_input[597], g_input[623]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[527]));
    dotproduct5 operation_conv528(.clk (clk), .rst (rst), .g_input ({g_input[568], g_input[569], g_input[596], g_input[598], g_input[624]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[528]));
    dotproduct5 operation_conv529(.clk (clk), .rst (rst), .g_input ({g_input[569], g_input[570], g_input[597], g_input[599], g_input[625]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[529]));
    dotproduct5 operation_conv530(.clk (clk), .rst (rst), .g_input ({g_input[570], g_input[571], g_input[598], g_input[600], g_input[626]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[530]));
    dotproduct5 operation_conv531(.clk (clk), .rst (rst), .g_input ({g_input[571], g_input[572], g_input[599], g_input[601], g_input[627]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[531]));
    dotproduct5 operation_conv532(.clk (clk), .rst (rst), .g_input ({g_input[572], g_input[573], g_input[600], g_input[602], g_input[628]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[532]));
    dotproduct5 operation_conv533(.clk (clk), .rst (rst), .g_input ({g_input[573], g_input[574], g_input[601], g_input[603], g_input[629]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[533]));
    dotproduct5 operation_conv534(.clk (clk), .rst (rst), .g_input ({g_input[574], g_input[575], g_input[602], g_input[604], g_input[630]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[534]));
    dotproduct5 operation_conv535(.clk (clk), .rst (rst), .g_input ({g_input[575], g_input[576], g_input[603], g_input[605], g_input[631]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[535]));
    dotproduct5 operation_conv536(.clk (clk), .rst (rst), .g_input ({g_input[576], g_input[577], g_input[604], g_input[606], g_input[632]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[536]));
    dotproduct5 operation_conv537(.clk (clk), .rst (rst), .g_input ({g_input[577], g_input[578], g_input[605], g_input[607], g_input[633]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[537]));
    dotproduct5 operation_conv538(.clk (clk), .rst (rst), .g_input ({g_input[578], g_input[579], g_input[606], g_input[608], g_input[634]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[538]));
    dotproduct5 operation_conv539(.clk (clk), .rst (rst), .g_input ({g_input[579], g_input[580], g_input[607], g_input[609], g_input[635]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[539]));
    dotproduct5 operation_conv540(.clk (clk), .rst (rst), .g_input ({g_input[580], g_input[581], g_input[608], g_input[610], g_input[636]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[540]));
    dotproduct5 operation_conv541(.clk (clk), .rst (rst), .g_input ({g_input[581], g_input[582], g_input[609], g_input[611], g_input[637]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[541]));
    dotproduct5 operation_conv542(.clk (clk), .rst (rst), .g_input ({g_input[582], g_input[583], g_input[610], g_input[612], g_input[638]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[542]));
    dotproduct5 operation_conv543(.clk (clk), .rst (rst), .g_input ({g_input[583], g_input[584], g_input[611], g_input[613], g_input[639]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[543]));
    dotproduct5 operation_conv544(.clk (clk), .rst (rst), .g_input ({g_input[584], g_input[585], g_input[612], g_input[614], g_input[640]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[544]));
    dotproduct5 operation_conv545(.clk (clk), .rst (rst), .g_input ({g_input[585], g_input[586], g_input[613], g_input[615], g_input[641]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[545]));
    dotproduct5 operation_conv546(.clk (clk), .rst (rst), .g_input ({g_input[588], g_input[589], g_input[616], g_input[618], g_input[644]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[546]));
    dotproduct5 operation_conv547(.clk (clk), .rst (rst), .g_input ({g_input[589], g_input[590], g_input[617], g_input[619], g_input[645]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[547]));
    dotproduct5 operation_conv548(.clk (clk), .rst (rst), .g_input ({g_input[590], g_input[591], g_input[618], g_input[620], g_input[646]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[548]));
    dotproduct5 operation_conv549(.clk (clk), .rst (rst), .g_input ({g_input[591], g_input[592], g_input[619], g_input[621], g_input[647]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[549]));
    dotproduct5 operation_conv550(.clk (clk), .rst (rst), .g_input ({g_input[592], g_input[593], g_input[620], g_input[622], g_input[648]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[550]));
    dotproduct5 operation_conv551(.clk (clk), .rst (rst), .g_input ({g_input[593], g_input[594], g_input[621], g_input[623], g_input[649]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[551]));
    dotproduct5 operation_conv552(.clk (clk), .rst (rst), .g_input ({g_input[594], g_input[595], g_input[622], g_input[624], g_input[650]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[552]));
    dotproduct5 operation_conv553(.clk (clk), .rst (rst), .g_input ({g_input[595], g_input[596], g_input[623], g_input[625], g_input[651]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[553]));
    dotproduct5 operation_conv554(.clk (clk), .rst (rst), .g_input ({g_input[596], g_input[597], g_input[624], g_input[626], g_input[652]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[554]));
    dotproduct5 operation_conv555(.clk (clk), .rst (rst), .g_input ({g_input[597], g_input[598], g_input[625], g_input[627], g_input[653]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[555]));
    dotproduct5 operation_conv556(.clk (clk), .rst (rst), .g_input ({g_input[598], g_input[599], g_input[626], g_input[628], g_input[654]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[556]));
    dotproduct5 operation_conv557(.clk (clk), .rst (rst), .g_input ({g_input[599], g_input[600], g_input[627], g_input[629], g_input[655]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[557]));
    dotproduct5 operation_conv558(.clk (clk), .rst (rst), .g_input ({g_input[600], g_input[601], g_input[628], g_input[630], g_input[656]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[558]));
    dotproduct5 operation_conv559(.clk (clk), .rst (rst), .g_input ({g_input[601], g_input[602], g_input[629], g_input[631], g_input[657]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[559]));
    dotproduct5 operation_conv560(.clk (clk), .rst (rst), .g_input ({g_input[602], g_input[603], g_input[630], g_input[632], g_input[658]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[560]));
    dotproduct5 operation_conv561(.clk (clk), .rst (rst), .g_input ({g_input[603], g_input[604], g_input[631], g_input[633], g_input[659]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[561]));
    dotproduct5 operation_conv562(.clk (clk), .rst (rst), .g_input ({g_input[604], g_input[605], g_input[632], g_input[634], g_input[660]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[562]));
    dotproduct5 operation_conv563(.clk (clk), .rst (rst), .g_input ({g_input[605], g_input[606], g_input[633], g_input[635], g_input[661]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[563]));
    dotproduct5 operation_conv564(.clk (clk), .rst (rst), .g_input ({g_input[606], g_input[607], g_input[634], g_input[636], g_input[662]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[564]));
    dotproduct5 operation_conv565(.clk (clk), .rst (rst), .g_input ({g_input[607], g_input[608], g_input[635], g_input[637], g_input[663]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[565]));
    dotproduct5 operation_conv566(.clk (clk), .rst (rst), .g_input ({g_input[608], g_input[609], g_input[636], g_input[638], g_input[664]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[566]));
    dotproduct5 operation_conv567(.clk (clk), .rst (rst), .g_input ({g_input[609], g_input[610], g_input[637], g_input[639], g_input[665]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[567]));
    dotproduct5 operation_conv568(.clk (clk), .rst (rst), .g_input ({g_input[610], g_input[611], g_input[638], g_input[640], g_input[666]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[568]));
    dotproduct5 operation_conv569(.clk (clk), .rst (rst), .g_input ({g_input[611], g_input[612], g_input[639], g_input[641], g_input[667]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[569]));
    dotproduct5 operation_conv570(.clk (clk), .rst (rst), .g_input ({g_input[612], g_input[613], g_input[640], g_input[642], g_input[668]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[570]));
    dotproduct5 operation_conv571(.clk (clk), .rst (rst), .g_input ({g_input[613], g_input[614], g_input[641], g_input[643], g_input[669]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[571]));
    dotproduct5 operation_conv572(.clk (clk), .rst (rst), .g_input ({g_input[616], g_input[617], g_input[644], g_input[646], g_input[672]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[572]));
    dotproduct5 operation_conv573(.clk (clk), .rst (rst), .g_input ({g_input[617], g_input[618], g_input[645], g_input[647], g_input[673]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[573]));
    dotproduct5 operation_conv574(.clk (clk), .rst (rst), .g_input ({g_input[618], g_input[619], g_input[646], g_input[648], g_input[674]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[574]));
    dotproduct5 operation_conv575(.clk (clk), .rst (rst), .g_input ({g_input[619], g_input[620], g_input[647], g_input[649], g_input[675]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[575]));
    dotproduct5 operation_conv576(.clk (clk), .rst (rst), .g_input ({g_input[620], g_input[621], g_input[648], g_input[650], g_input[676]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[576]));
    dotproduct5 operation_conv577(.clk (clk), .rst (rst), .g_input ({g_input[621], g_input[622], g_input[649], g_input[651], g_input[677]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[577]));
    dotproduct5 operation_conv578(.clk (clk), .rst (rst), .g_input ({g_input[622], g_input[623], g_input[650], g_input[652], g_input[678]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[578]));
    dotproduct5 operation_conv579(.clk (clk), .rst (rst), .g_input ({g_input[623], g_input[624], g_input[651], g_input[653], g_input[679]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[579]));
    dotproduct5 operation_conv580(.clk (clk), .rst (rst), .g_input ({g_input[624], g_input[625], g_input[652], g_input[654], g_input[680]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[580]));
    dotproduct5 operation_conv581(.clk (clk), .rst (rst), .g_input ({g_input[625], g_input[626], g_input[653], g_input[655], g_input[681]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[581]));
    dotproduct5 operation_conv582(.clk (clk), .rst (rst), .g_input ({g_input[626], g_input[627], g_input[654], g_input[656], g_input[682]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[582]));
    dotproduct5 operation_conv583(.clk (clk), .rst (rst), .g_input ({g_input[627], g_input[628], g_input[655], g_input[657], g_input[683]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[583]));
    dotproduct5 operation_conv584(.clk (clk), .rst (rst), .g_input ({g_input[628], g_input[629], g_input[656], g_input[658], g_input[684]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[584]));
    dotproduct5 operation_conv585(.clk (clk), .rst (rst), .g_input ({g_input[629], g_input[630], g_input[657], g_input[659], g_input[685]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[585]));
    dotproduct5 operation_conv586(.clk (clk), .rst (rst), .g_input ({g_input[630], g_input[631], g_input[658], g_input[660], g_input[686]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[586]));
    dotproduct5 operation_conv587(.clk (clk), .rst (rst), .g_input ({g_input[631], g_input[632], g_input[659], g_input[661], g_input[687]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[587]));
    dotproduct5 operation_conv588(.clk (clk), .rst (rst), .g_input ({g_input[632], g_input[633], g_input[660], g_input[662], g_input[688]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[588]));
    dotproduct5 operation_conv589(.clk (clk), .rst (rst), .g_input ({g_input[633], g_input[634], g_input[661], g_input[663], g_input[689]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[589]));
    dotproduct5 operation_conv590(.clk (clk), .rst (rst), .g_input ({g_input[634], g_input[635], g_input[662], g_input[664], g_input[690]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[590]));
    dotproduct5 operation_conv591(.clk (clk), .rst (rst), .g_input ({g_input[635], g_input[636], g_input[663], g_input[665], g_input[691]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[591]));
    dotproduct5 operation_conv592(.clk (clk), .rst (rst), .g_input ({g_input[636], g_input[637], g_input[664], g_input[666], g_input[692]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[592]));
    dotproduct5 operation_conv593(.clk (clk), .rst (rst), .g_input ({g_input[637], g_input[638], g_input[665], g_input[667], g_input[693]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[593]));
    dotproduct5 operation_conv594(.clk (clk), .rst (rst), .g_input ({g_input[638], g_input[639], g_input[666], g_input[668], g_input[694]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[594]));
    dotproduct5 operation_conv595(.clk (clk), .rst (rst), .g_input ({g_input[639], g_input[640], g_input[667], g_input[669], g_input[695]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[595]));
    dotproduct5 operation_conv596(.clk (clk), .rst (rst), .g_input ({g_input[640], g_input[641], g_input[668], g_input[670], g_input[696]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[596]));
    dotproduct5 operation_conv597(.clk (clk), .rst (rst), .g_input ({g_input[641], g_input[642], g_input[669], g_input[671], g_input[697]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[597]));
    dotproduct5 operation_conv598(.clk (clk), .rst (rst), .g_input ({g_input[644], g_input[645], g_input[672], g_input[674], g_input[700]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[598]));
    dotproduct5 operation_conv599(.clk (clk), .rst (rst), .g_input ({g_input[645], g_input[646], g_input[673], g_input[675], g_input[701]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[599]));
    dotproduct5 operation_conv600(.clk (clk), .rst (rst), .g_input ({g_input[646], g_input[647], g_input[674], g_input[676], g_input[702]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[600]));
    dotproduct5 operation_conv601(.clk (clk), .rst (rst), .g_input ({g_input[647], g_input[648], g_input[675], g_input[677], g_input[703]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[601]));
    dotproduct5 operation_conv602(.clk (clk), .rst (rst), .g_input ({g_input[648], g_input[649], g_input[676], g_input[678], g_input[704]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[602]));
    dotproduct5 operation_conv603(.clk (clk), .rst (rst), .g_input ({g_input[649], g_input[650], g_input[677], g_input[679], g_input[705]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[603]));
    dotproduct5 operation_conv604(.clk (clk), .rst (rst), .g_input ({g_input[650], g_input[651], g_input[678], g_input[680], g_input[706]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[604]));
    dotproduct5 operation_conv605(.clk (clk), .rst (rst), .g_input ({g_input[651], g_input[652], g_input[679], g_input[681], g_input[707]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[605]));
    dotproduct5 operation_conv606(.clk (clk), .rst (rst), .g_input ({g_input[652], g_input[653], g_input[680], g_input[682], g_input[708]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[606]));
    dotproduct5 operation_conv607(.clk (clk), .rst (rst), .g_input ({g_input[653], g_input[654], g_input[681], g_input[683], g_input[709]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[607]));
    dotproduct5 operation_conv608(.clk (clk), .rst (rst), .g_input ({g_input[654], g_input[655], g_input[682], g_input[684], g_input[710]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[608]));
    dotproduct5 operation_conv609(.clk (clk), .rst (rst), .g_input ({g_input[655], g_input[656], g_input[683], g_input[685], g_input[711]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[609]));
    dotproduct5 operation_conv610(.clk (clk), .rst (rst), .g_input ({g_input[656], g_input[657], g_input[684], g_input[686], g_input[712]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[610]));
    dotproduct5 operation_conv611(.clk (clk), .rst (rst), .g_input ({g_input[657], g_input[658], g_input[685], g_input[687], g_input[713]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[611]));
    dotproduct5 operation_conv612(.clk (clk), .rst (rst), .g_input ({g_input[658], g_input[659], g_input[686], g_input[688], g_input[714]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[612]));
    dotproduct5 operation_conv613(.clk (clk), .rst (rst), .g_input ({g_input[659], g_input[660], g_input[687], g_input[689], g_input[715]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[613]));
    dotproduct5 operation_conv614(.clk (clk), .rst (rst), .g_input ({g_input[660], g_input[661], g_input[688], g_input[690], g_input[716]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[614]));
    dotproduct5 operation_conv615(.clk (clk), .rst (rst), .g_input ({g_input[661], g_input[662], g_input[689], g_input[691], g_input[717]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[615]));
    dotproduct5 operation_conv616(.clk (clk), .rst (rst), .g_input ({g_input[662], g_input[663], g_input[690], g_input[692], g_input[718]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[616]));
    dotproduct5 operation_conv617(.clk (clk), .rst (rst), .g_input ({g_input[663], g_input[664], g_input[691], g_input[693], g_input[719]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[617]));
    dotproduct5 operation_conv618(.clk (clk), .rst (rst), .g_input ({g_input[664], g_input[665], g_input[692], g_input[694], g_input[720]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[618]));
    dotproduct5 operation_conv619(.clk (clk), .rst (rst), .g_input ({g_input[665], g_input[666], g_input[693], g_input[695], g_input[721]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[619]));
    dotproduct5 operation_conv620(.clk (clk), .rst (rst), .g_input ({g_input[666], g_input[667], g_input[694], g_input[696], g_input[722]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[620]));
    dotproduct5 operation_conv621(.clk (clk), .rst (rst), .g_input ({g_input[667], g_input[668], g_input[695], g_input[697], g_input[723]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[621]));
    dotproduct5 operation_conv622(.clk (clk), .rst (rst), .g_input ({g_input[668], g_input[669], g_input[696], g_input[698], g_input[724]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[622]));
    dotproduct5 operation_conv623(.clk (clk), .rst (rst), .g_input ({g_input[669], g_input[670], g_input[697], g_input[699], g_input[725]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[623]));
    dotproduct5 operation_conv624(.clk (clk), .rst (rst), .g_input ({g_input[672], g_input[673], g_input[700], g_input[702], g_input[728]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[624]));
    dotproduct5 operation_conv625(.clk (clk), .rst (rst), .g_input ({g_input[673], g_input[674], g_input[701], g_input[703], g_input[729]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[625]));
    dotproduct5 operation_conv626(.clk (clk), .rst (rst), .g_input ({g_input[674], g_input[675], g_input[702], g_input[704], g_input[730]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[626]));
    dotproduct5 operation_conv627(.clk (clk), .rst (rst), .g_input ({g_input[675], g_input[676], g_input[703], g_input[705], g_input[731]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[627]));
    dotproduct5 operation_conv628(.clk (clk), .rst (rst), .g_input ({g_input[676], g_input[677], g_input[704], g_input[706], g_input[732]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[628]));
    dotproduct5 operation_conv629(.clk (clk), .rst (rst), .g_input ({g_input[677], g_input[678], g_input[705], g_input[707], g_input[733]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[629]));
    dotproduct5 operation_conv630(.clk (clk), .rst (rst), .g_input ({g_input[678], g_input[679], g_input[706], g_input[708], g_input[734]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[630]));
    dotproduct5 operation_conv631(.clk (clk), .rst (rst), .g_input ({g_input[679], g_input[680], g_input[707], g_input[709], g_input[735]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[631]));
    dotproduct5 operation_conv632(.clk (clk), .rst (rst), .g_input ({g_input[680], g_input[681], g_input[708], g_input[710], g_input[736]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[632]));
    dotproduct5 operation_conv633(.clk (clk), .rst (rst), .g_input ({g_input[681], g_input[682], g_input[709], g_input[711], g_input[737]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[633]));
    dotproduct5 operation_conv634(.clk (clk), .rst (rst), .g_input ({g_input[682], g_input[683], g_input[710], g_input[712], g_input[738]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[634]));
    dotproduct5 operation_conv635(.clk (clk), .rst (rst), .g_input ({g_input[683], g_input[684], g_input[711], g_input[713], g_input[739]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[635]));
    dotproduct5 operation_conv636(.clk (clk), .rst (rst), .g_input ({g_input[684], g_input[685], g_input[712], g_input[714], g_input[740]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[636]));
    dotproduct5 operation_conv637(.clk (clk), .rst (rst), .g_input ({g_input[685], g_input[686], g_input[713], g_input[715], g_input[741]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[637]));
    dotproduct5 operation_conv638(.clk (clk), .rst (rst), .g_input ({g_input[686], g_input[687], g_input[714], g_input[716], g_input[742]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[638]));
    dotproduct5 operation_conv639(.clk (clk), .rst (rst), .g_input ({g_input[687], g_input[688], g_input[715], g_input[717], g_input[743]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[639]));
    dotproduct5 operation_conv640(.clk (clk), .rst (rst), .g_input ({g_input[688], g_input[689], g_input[716], g_input[718], g_input[744]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[640]));
    dotproduct5 operation_conv641(.clk (clk), .rst (rst), .g_input ({g_input[689], g_input[690], g_input[717], g_input[719], g_input[745]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[641]));
    dotproduct5 operation_conv642(.clk (clk), .rst (rst), .g_input ({g_input[690], g_input[691], g_input[718], g_input[720], g_input[746]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[642]));
    dotproduct5 operation_conv643(.clk (clk), .rst (rst), .g_input ({g_input[691], g_input[692], g_input[719], g_input[721], g_input[747]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[643]));
    dotproduct5 operation_conv644(.clk (clk), .rst (rst), .g_input ({g_input[692], g_input[693], g_input[720], g_input[722], g_input[748]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[644]));
    dotproduct5 operation_conv645(.clk (clk), .rst (rst), .g_input ({g_input[693], g_input[694], g_input[721], g_input[723], g_input[749]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[645]));
    dotproduct5 operation_conv646(.clk (clk), .rst (rst), .g_input ({g_input[694], g_input[695], g_input[722], g_input[724], g_input[750]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[646]));
    dotproduct5 operation_conv647(.clk (clk), .rst (rst), .g_input ({g_input[695], g_input[696], g_input[723], g_input[725], g_input[751]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[647]));
    dotproduct5 operation_conv648(.clk (clk), .rst (rst), .g_input ({g_input[696], g_input[697], g_input[724], g_input[726], g_input[752]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[648]));
    dotproduct5 operation_conv649(.clk (clk), .rst (rst), .g_input ({g_input[697], g_input[698], g_input[725], g_input[727], g_input[753]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[649]));
    dotproduct5 operation_conv650(.clk (clk), .rst (rst), .g_input ({g_input[700], g_input[701], g_input[728], g_input[730], g_input[756]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[650]));
    dotproduct5 operation_conv651(.clk (clk), .rst (rst), .g_input ({g_input[701], g_input[702], g_input[729], g_input[731], g_input[757]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[651]));
    dotproduct5 operation_conv652(.clk (clk), .rst (rst), .g_input ({g_input[702], g_input[703], g_input[730], g_input[732], g_input[758]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[652]));
    dotproduct5 operation_conv653(.clk (clk), .rst (rst), .g_input ({g_input[703], g_input[704], g_input[731], g_input[733], g_input[759]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[653]));
    dotproduct5 operation_conv654(.clk (clk), .rst (rst), .g_input ({g_input[704], g_input[705], g_input[732], g_input[734], g_input[760]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[654]));
    dotproduct5 operation_conv655(.clk (clk), .rst (rst), .g_input ({g_input[705], g_input[706], g_input[733], g_input[735], g_input[761]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[655]));
    dotproduct5 operation_conv656(.clk (clk), .rst (rst), .g_input ({g_input[706], g_input[707], g_input[734], g_input[736], g_input[762]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[656]));
    dotproduct5 operation_conv657(.clk (clk), .rst (rst), .g_input ({g_input[707], g_input[708], g_input[735], g_input[737], g_input[763]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[657]));
    dotproduct5 operation_conv658(.clk (clk), .rst (rst), .g_input ({g_input[708], g_input[709], g_input[736], g_input[738], g_input[764]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[658]));
    dotproduct5 operation_conv659(.clk (clk), .rst (rst), .g_input ({g_input[709], g_input[710], g_input[737], g_input[739], g_input[765]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[659]));
    dotproduct5 operation_conv660(.clk (clk), .rst (rst), .g_input ({g_input[710], g_input[711], g_input[738], g_input[740], g_input[766]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[660]));
    dotproduct5 operation_conv661(.clk (clk), .rst (rst), .g_input ({g_input[711], g_input[712], g_input[739], g_input[741], g_input[767]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[661]));
    dotproduct5 operation_conv662(.clk (clk), .rst (rst), .g_input ({g_input[712], g_input[713], g_input[740], g_input[742], g_input[768]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[662]));
    dotproduct5 operation_conv663(.clk (clk), .rst (rst), .g_input ({g_input[713], g_input[714], g_input[741], g_input[743], g_input[769]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[663]));
    dotproduct5 operation_conv664(.clk (clk), .rst (rst), .g_input ({g_input[714], g_input[715], g_input[742], g_input[744], g_input[770]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[664]));
    dotproduct5 operation_conv665(.clk (clk), .rst (rst), .g_input ({g_input[715], g_input[716], g_input[743], g_input[745], g_input[771]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[665]));
    dotproduct5 operation_conv666(.clk (clk), .rst (rst), .g_input ({g_input[716], g_input[717], g_input[744], g_input[746], g_input[772]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[666]));
    dotproduct5 operation_conv667(.clk (clk), .rst (rst), .g_input ({g_input[717], g_input[718], g_input[745], g_input[747], g_input[773]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[667]));
    dotproduct5 operation_conv668(.clk (clk), .rst (rst), .g_input ({g_input[718], g_input[719], g_input[746], g_input[748], g_input[774]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[668]));
    dotproduct5 operation_conv669(.clk (clk), .rst (rst), .g_input ({g_input[719], g_input[720], g_input[747], g_input[749], g_input[775]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[669]));
    dotproduct5 operation_conv670(.clk (clk), .rst (rst), .g_input ({g_input[720], g_input[721], g_input[748], g_input[750], g_input[776]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[670]));
    dotproduct5 operation_conv671(.clk (clk), .rst (rst), .g_input ({g_input[721], g_input[722], g_input[749], g_input[751], g_input[777]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[671]));
    dotproduct5 operation_conv672(.clk (clk), .rst (rst), .g_input ({g_input[722], g_input[723], g_input[750], g_input[752], g_input[778]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[672]));
    dotproduct5 operation_conv673(.clk (clk), .rst (rst), .g_input ({g_input[723], g_input[724], g_input[751], g_input[753], g_input[779]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[673]));
    dotproduct5 operation_conv674(.clk (clk), .rst (rst), .g_input ({g_input[724], g_input[725], g_input[752], g_input[754], g_input[780]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[674]));
    dotproduct5 operation_conv675(.clk (clk), .rst (rst), .g_input ({g_input[725], g_input[726], g_input[753], g_input[755], g_input[781]}), .e_input({e_input[0], e_input[1], e_input[3], e_input[5], e_input[6]}), .o (conv1_0_0[675]));
    assign conv1_res = {conv1_0_0};


        maxpool1 operation_mp1676(
            .clk   (clk),
            .rst   (rst),
            .g_input (conv1_res[675:0]),
            .e_input (1'b0),
            .o     (mp1_0)
        );
        assign mp1_res = {mp1_0};

    dotproduct15 operation_conv677(.clk (clk), .rst (rst), .g_input ({mp1_res[0], mp1_res[1], mp1_res[2], mp1_res[3], mp1_res[14], mp1_res[15], mp1_res[17], mp1_res[28], mp1_res[29], mp1_res[39], mp1_res[40], mp1_res[41], mp1_res[52], mp1_res[54], mp1_res[56]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[0]));
    dotproduct15 operation_conv678(.clk (clk), .rst (rst), .g_input ({mp1_res[1], mp1_res[2], mp1_res[3], mp1_res[4], mp1_res[15], mp1_res[16], mp1_res[18], mp1_res[29], mp1_res[30], mp1_res[40], mp1_res[41], mp1_res[42], mp1_res[53], mp1_res[55], mp1_res[57]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[1]));
    dotproduct15 operation_conv679(.clk (clk), .rst (rst), .g_input ({mp1_res[2], mp1_res[3], mp1_res[4], mp1_res[5], mp1_res[16], mp1_res[17], mp1_res[19], mp1_res[30], mp1_res[31], mp1_res[41], mp1_res[42], mp1_res[43], mp1_res[54], mp1_res[56], mp1_res[58]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[2]));
    dotproduct15 operation_conv680(.clk (clk), .rst (rst), .g_input ({mp1_res[3], mp1_res[4], mp1_res[5], mp1_res[6], mp1_res[17], mp1_res[18], mp1_res[20], mp1_res[31], mp1_res[32], mp1_res[42], mp1_res[43], mp1_res[44], mp1_res[55], mp1_res[57], mp1_res[59]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[3]));
    dotproduct15 operation_conv681(.clk (clk), .rst (rst), .g_input ({mp1_res[4], mp1_res[5], mp1_res[6], mp1_res[7], mp1_res[18], mp1_res[19], mp1_res[21], mp1_res[32], mp1_res[33], mp1_res[43], mp1_res[44], mp1_res[45], mp1_res[56], mp1_res[58], mp1_res[60]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[4]));
    dotproduct15 operation_conv682(.clk (clk), .rst (rst), .g_input ({mp1_res[5], mp1_res[6], mp1_res[7], mp1_res[8], mp1_res[19], mp1_res[20], mp1_res[22], mp1_res[33], mp1_res[34], mp1_res[44], mp1_res[45], mp1_res[46], mp1_res[57], mp1_res[59], mp1_res[61]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[5]));
    dotproduct15 operation_conv683(.clk (clk), .rst (rst), .g_input ({mp1_res[6], mp1_res[7], mp1_res[8], mp1_res[9], mp1_res[20], mp1_res[21], mp1_res[23], mp1_res[34], mp1_res[35], mp1_res[45], mp1_res[46], mp1_res[47], mp1_res[58], mp1_res[60], mp1_res[62]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[6]));
    dotproduct15 operation_conv684(.clk (clk), .rst (rst), .g_input ({mp1_res[7], mp1_res[8], mp1_res[9], mp1_res[10], mp1_res[21], mp1_res[22], mp1_res[24], mp1_res[35], mp1_res[36], mp1_res[46], mp1_res[47], mp1_res[48], mp1_res[59], mp1_res[61], mp1_res[63]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[7]));
    dotproduct15 operation_conv685(.clk (clk), .rst (rst), .g_input ({mp1_res[8], mp1_res[9], mp1_res[10], mp1_res[11], mp1_res[22], mp1_res[23], mp1_res[25], mp1_res[36], mp1_res[37], mp1_res[47], mp1_res[48], mp1_res[49], mp1_res[60], mp1_res[62], mp1_res[64]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[8]));
    dotproduct15 operation_conv686(.clk (clk), .rst (rst), .g_input ({mp1_res[13], mp1_res[14], mp1_res[15], mp1_res[16], mp1_res[27], mp1_res[28], mp1_res[30], mp1_res[41], mp1_res[42], mp1_res[52], mp1_res[53], mp1_res[54], mp1_res[65], mp1_res[67], mp1_res[69]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[9]));
    dotproduct15 operation_conv687(.clk (clk), .rst (rst), .g_input ({mp1_res[14], mp1_res[15], mp1_res[16], mp1_res[17], mp1_res[28], mp1_res[29], mp1_res[31], mp1_res[42], mp1_res[43], mp1_res[53], mp1_res[54], mp1_res[55], mp1_res[66], mp1_res[68], mp1_res[70]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[10]));
    dotproduct15 operation_conv688(.clk (clk), .rst (rst), .g_input ({mp1_res[15], mp1_res[16], mp1_res[17], mp1_res[18], mp1_res[29], mp1_res[30], mp1_res[32], mp1_res[43], mp1_res[44], mp1_res[54], mp1_res[55], mp1_res[56], mp1_res[67], mp1_res[69], mp1_res[71]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[11]));
    dotproduct15 operation_conv689(.clk (clk), .rst (rst), .g_input ({mp1_res[16], mp1_res[17], mp1_res[18], mp1_res[19], mp1_res[30], mp1_res[31], mp1_res[33], mp1_res[44], mp1_res[45], mp1_res[55], mp1_res[56], mp1_res[57], mp1_res[68], mp1_res[70], mp1_res[72]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[12]));
    dotproduct15 operation_conv690(.clk (clk), .rst (rst), .g_input ({mp1_res[17], mp1_res[18], mp1_res[19], mp1_res[20], mp1_res[31], mp1_res[32], mp1_res[34], mp1_res[45], mp1_res[46], mp1_res[56], mp1_res[57], mp1_res[58], mp1_res[69], mp1_res[71], mp1_res[73]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[13]));
    dotproduct15 operation_conv691(.clk (clk), .rst (rst), .g_input ({mp1_res[18], mp1_res[19], mp1_res[20], mp1_res[21], mp1_res[32], mp1_res[33], mp1_res[35], mp1_res[46], mp1_res[47], mp1_res[57], mp1_res[58], mp1_res[59], mp1_res[70], mp1_res[72], mp1_res[74]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[14]));
    dotproduct15 operation_conv692(.clk (clk), .rst (rst), .g_input ({mp1_res[19], mp1_res[20], mp1_res[21], mp1_res[22], mp1_res[33], mp1_res[34], mp1_res[36], mp1_res[47], mp1_res[48], mp1_res[58], mp1_res[59], mp1_res[60], mp1_res[71], mp1_res[73], mp1_res[75]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[15]));
    dotproduct15 operation_conv693(.clk (clk), .rst (rst), .g_input ({mp1_res[20], mp1_res[21], mp1_res[22], mp1_res[23], mp1_res[34], mp1_res[35], mp1_res[37], mp1_res[48], mp1_res[49], mp1_res[59], mp1_res[60], mp1_res[61], mp1_res[72], mp1_res[74], mp1_res[76]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[16]));
    dotproduct15 operation_conv694(.clk (clk), .rst (rst), .g_input ({mp1_res[21], mp1_res[22], mp1_res[23], mp1_res[24], mp1_res[35], mp1_res[36], mp1_res[38], mp1_res[49], mp1_res[50], mp1_res[60], mp1_res[61], mp1_res[62], mp1_res[73], mp1_res[75], mp1_res[77]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[17]));
    dotproduct15 operation_conv695(.clk (clk), .rst (rst), .g_input ({mp1_res[26], mp1_res[27], mp1_res[28], mp1_res[29], mp1_res[40], mp1_res[41], mp1_res[43], mp1_res[54], mp1_res[55], mp1_res[65], mp1_res[66], mp1_res[67], mp1_res[78], mp1_res[80], mp1_res[82]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[18]));
    dotproduct15 operation_conv696(.clk (clk), .rst (rst), .g_input ({mp1_res[27], mp1_res[28], mp1_res[29], mp1_res[30], mp1_res[41], mp1_res[42], mp1_res[44], mp1_res[55], mp1_res[56], mp1_res[66], mp1_res[67], mp1_res[68], mp1_res[79], mp1_res[81], mp1_res[83]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[19]));
    dotproduct15 operation_conv697(.clk (clk), .rst (rst), .g_input ({mp1_res[28], mp1_res[29], mp1_res[30], mp1_res[31], mp1_res[42], mp1_res[43], mp1_res[45], mp1_res[56], mp1_res[57], mp1_res[67], mp1_res[68], mp1_res[69], mp1_res[80], mp1_res[82], mp1_res[84]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[20]));
    dotproduct15 operation_conv698(.clk (clk), .rst (rst), .g_input ({mp1_res[29], mp1_res[30], mp1_res[31], mp1_res[32], mp1_res[43], mp1_res[44], mp1_res[46], mp1_res[57], mp1_res[58], mp1_res[68], mp1_res[69], mp1_res[70], mp1_res[81], mp1_res[83], mp1_res[85]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[21]));
    dotproduct15 operation_conv699(.clk (clk), .rst (rst), .g_input ({mp1_res[30], mp1_res[31], mp1_res[32], mp1_res[33], mp1_res[44], mp1_res[45], mp1_res[47], mp1_res[58], mp1_res[59], mp1_res[69], mp1_res[70], mp1_res[71], mp1_res[82], mp1_res[84], mp1_res[86]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[22]));
    dotproduct15 operation_conv700(.clk (clk), .rst (rst), .g_input ({mp1_res[31], mp1_res[32], mp1_res[33], mp1_res[34], mp1_res[45], mp1_res[46], mp1_res[48], mp1_res[59], mp1_res[60], mp1_res[70], mp1_res[71], mp1_res[72], mp1_res[83], mp1_res[85], mp1_res[87]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[23]));
    dotproduct15 operation_conv701(.clk (clk), .rst (rst), .g_input ({mp1_res[32], mp1_res[33], mp1_res[34], mp1_res[35], mp1_res[46], mp1_res[47], mp1_res[49], mp1_res[60], mp1_res[61], mp1_res[71], mp1_res[72], mp1_res[73], mp1_res[84], mp1_res[86], mp1_res[88]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[24]));
    dotproduct15 operation_conv702(.clk (clk), .rst (rst), .g_input ({mp1_res[33], mp1_res[34], mp1_res[35], mp1_res[36], mp1_res[47], mp1_res[48], mp1_res[50], mp1_res[61], mp1_res[62], mp1_res[72], mp1_res[73], mp1_res[74], mp1_res[85], mp1_res[87], mp1_res[89]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[25]));
    dotproduct15 operation_conv703(.clk (clk), .rst (rst), .g_input ({mp1_res[34], mp1_res[35], mp1_res[36], mp1_res[37], mp1_res[48], mp1_res[49], mp1_res[51], mp1_res[62], mp1_res[63], mp1_res[73], mp1_res[74], mp1_res[75], mp1_res[86], mp1_res[88], mp1_res[90]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[26]));
    dotproduct15 operation_conv704(.clk (clk), .rst (rst), .g_input ({mp1_res[39], mp1_res[40], mp1_res[41], mp1_res[42], mp1_res[53], mp1_res[54], mp1_res[56], mp1_res[67], mp1_res[68], mp1_res[78], mp1_res[79], mp1_res[80], mp1_res[91], mp1_res[93], mp1_res[95]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[27]));
    dotproduct15 operation_conv705(.clk (clk), .rst (rst), .g_input ({mp1_res[40], mp1_res[41], mp1_res[42], mp1_res[43], mp1_res[54], mp1_res[55], mp1_res[57], mp1_res[68], mp1_res[69], mp1_res[79], mp1_res[80], mp1_res[81], mp1_res[92], mp1_res[94], mp1_res[96]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[28]));
    dotproduct15 operation_conv706(.clk (clk), .rst (rst), .g_input ({mp1_res[41], mp1_res[42], mp1_res[43], mp1_res[44], mp1_res[55], mp1_res[56], mp1_res[58], mp1_res[69], mp1_res[70], mp1_res[80], mp1_res[81], mp1_res[82], mp1_res[93], mp1_res[95], mp1_res[97]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[29]));
    dotproduct15 operation_conv707(.clk (clk), .rst (rst), .g_input ({mp1_res[42], mp1_res[43], mp1_res[44], mp1_res[45], mp1_res[56], mp1_res[57], mp1_res[59], mp1_res[70], mp1_res[71], mp1_res[81], mp1_res[82], mp1_res[83], mp1_res[94], mp1_res[96], mp1_res[98]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[30]));
    dotproduct15 operation_conv708(.clk (clk), .rst (rst), .g_input ({mp1_res[43], mp1_res[44], mp1_res[45], mp1_res[46], mp1_res[57], mp1_res[58], mp1_res[60], mp1_res[71], mp1_res[72], mp1_res[82], mp1_res[83], mp1_res[84], mp1_res[95], mp1_res[97], mp1_res[99]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[31]));
    dotproduct15 operation_conv709(.clk (clk), .rst (rst), .g_input ({mp1_res[44], mp1_res[45], mp1_res[46], mp1_res[47], mp1_res[58], mp1_res[59], mp1_res[61], mp1_res[72], mp1_res[73], mp1_res[83], mp1_res[84], mp1_res[85], mp1_res[96], mp1_res[98], mp1_res[100]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[32]));
    dotproduct15 operation_conv710(.clk (clk), .rst (rst), .g_input ({mp1_res[45], mp1_res[46], mp1_res[47], mp1_res[48], mp1_res[59], mp1_res[60], mp1_res[62], mp1_res[73], mp1_res[74], mp1_res[84], mp1_res[85], mp1_res[86], mp1_res[97], mp1_res[99], mp1_res[101]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[33]));
    dotproduct15 operation_conv711(.clk (clk), .rst (rst), .g_input ({mp1_res[46], mp1_res[47], mp1_res[48], mp1_res[49], mp1_res[60], mp1_res[61], mp1_res[63], mp1_res[74], mp1_res[75], mp1_res[85], mp1_res[86], mp1_res[87], mp1_res[98], mp1_res[100], mp1_res[102]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[34]));
    dotproduct15 operation_conv712(.clk (clk), .rst (rst), .g_input ({mp1_res[47], mp1_res[48], mp1_res[49], mp1_res[50], mp1_res[61], mp1_res[62], mp1_res[64], mp1_res[75], mp1_res[76], mp1_res[86], mp1_res[87], mp1_res[88], mp1_res[99], mp1_res[101], mp1_res[103]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[35]));
    dotproduct15 operation_conv713(.clk (clk), .rst (rst), .g_input ({mp1_res[52], mp1_res[53], mp1_res[54], mp1_res[55], mp1_res[66], mp1_res[67], mp1_res[69], mp1_res[80], mp1_res[81], mp1_res[91], mp1_res[92], mp1_res[93], mp1_res[104], mp1_res[106], mp1_res[108]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[36]));
    dotproduct15 operation_conv714(.clk (clk), .rst (rst), .g_input ({mp1_res[53], mp1_res[54], mp1_res[55], mp1_res[56], mp1_res[67], mp1_res[68], mp1_res[70], mp1_res[81], mp1_res[82], mp1_res[92], mp1_res[93], mp1_res[94], mp1_res[105], mp1_res[107], mp1_res[109]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[37]));
    dotproduct15 operation_conv715(.clk (clk), .rst (rst), .g_input ({mp1_res[54], mp1_res[55], mp1_res[56], mp1_res[57], mp1_res[68], mp1_res[69], mp1_res[71], mp1_res[82], mp1_res[83], mp1_res[93], mp1_res[94], mp1_res[95], mp1_res[106], mp1_res[108], mp1_res[110]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[38]));
    dotproduct15 operation_conv716(.clk (clk), .rst (rst), .g_input ({mp1_res[55], mp1_res[56], mp1_res[57], mp1_res[58], mp1_res[69], mp1_res[70], mp1_res[72], mp1_res[83], mp1_res[84], mp1_res[94], mp1_res[95], mp1_res[96], mp1_res[107], mp1_res[109], mp1_res[111]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[39]));
    dotproduct15 operation_conv717(.clk (clk), .rst (rst), .g_input ({mp1_res[56], mp1_res[57], mp1_res[58], mp1_res[59], mp1_res[70], mp1_res[71], mp1_res[73], mp1_res[84], mp1_res[85], mp1_res[95], mp1_res[96], mp1_res[97], mp1_res[108], mp1_res[110], mp1_res[112]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[40]));
    dotproduct15 operation_conv718(.clk (clk), .rst (rst), .g_input ({mp1_res[57], mp1_res[58], mp1_res[59], mp1_res[60], mp1_res[71], mp1_res[72], mp1_res[74], mp1_res[85], mp1_res[86], mp1_res[96], mp1_res[97], mp1_res[98], mp1_res[109], mp1_res[111], mp1_res[113]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[41]));
    dotproduct15 operation_conv719(.clk (clk), .rst (rst), .g_input ({mp1_res[58], mp1_res[59], mp1_res[60], mp1_res[61], mp1_res[72], mp1_res[73], mp1_res[75], mp1_res[86], mp1_res[87], mp1_res[97], mp1_res[98], mp1_res[99], mp1_res[110], mp1_res[112], mp1_res[114]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[42]));
    dotproduct15 operation_conv720(.clk (clk), .rst (rst), .g_input ({mp1_res[59], mp1_res[60], mp1_res[61], mp1_res[62], mp1_res[73], mp1_res[74], mp1_res[76], mp1_res[87], mp1_res[88], mp1_res[98], mp1_res[99], mp1_res[100], mp1_res[111], mp1_res[113], mp1_res[115]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[43]));
    dotproduct15 operation_conv721(.clk (clk), .rst (rst), .g_input ({mp1_res[60], mp1_res[61], mp1_res[62], mp1_res[63], mp1_res[74], mp1_res[75], mp1_res[77], mp1_res[88], mp1_res[89], mp1_res[99], mp1_res[100], mp1_res[101], mp1_res[112], mp1_res[114], mp1_res[116]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[44]));
    dotproduct15 operation_conv722(.clk (clk), .rst (rst), .g_input ({mp1_res[65], mp1_res[66], mp1_res[67], mp1_res[68], mp1_res[79], mp1_res[80], mp1_res[82], mp1_res[93], mp1_res[94], mp1_res[104], mp1_res[105], mp1_res[106], mp1_res[117], mp1_res[119], mp1_res[121]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[45]));
    dotproduct15 operation_conv723(.clk (clk), .rst (rst), .g_input ({mp1_res[66], mp1_res[67], mp1_res[68], mp1_res[69], mp1_res[80], mp1_res[81], mp1_res[83], mp1_res[94], mp1_res[95], mp1_res[105], mp1_res[106], mp1_res[107], mp1_res[118], mp1_res[120], mp1_res[122]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[46]));
    dotproduct15 operation_conv724(.clk (clk), .rst (rst), .g_input ({mp1_res[67], mp1_res[68], mp1_res[69], mp1_res[70], mp1_res[81], mp1_res[82], mp1_res[84], mp1_res[95], mp1_res[96], mp1_res[106], mp1_res[107], mp1_res[108], mp1_res[119], mp1_res[121], mp1_res[123]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[47]));
    dotproduct15 operation_conv725(.clk (clk), .rst (rst), .g_input ({mp1_res[68], mp1_res[69], mp1_res[70], mp1_res[71], mp1_res[82], mp1_res[83], mp1_res[85], mp1_res[96], mp1_res[97], mp1_res[107], mp1_res[108], mp1_res[109], mp1_res[120], mp1_res[122], mp1_res[124]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[48]));
    dotproduct15 operation_conv726(.clk (clk), .rst (rst), .g_input ({mp1_res[69], mp1_res[70], mp1_res[71], mp1_res[72], mp1_res[83], mp1_res[84], mp1_res[86], mp1_res[97], mp1_res[98], mp1_res[108], mp1_res[109], mp1_res[110], mp1_res[121], mp1_res[123], mp1_res[125]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[49]));
    dotproduct15 operation_conv727(.clk (clk), .rst (rst), .g_input ({mp1_res[70], mp1_res[71], mp1_res[72], mp1_res[73], mp1_res[84], mp1_res[85], mp1_res[87], mp1_res[98], mp1_res[99], mp1_res[109], mp1_res[110], mp1_res[111], mp1_res[122], mp1_res[124], mp1_res[126]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[50]));
    dotproduct15 operation_conv728(.clk (clk), .rst (rst), .g_input ({mp1_res[71], mp1_res[72], mp1_res[73], mp1_res[74], mp1_res[85], mp1_res[86], mp1_res[88], mp1_res[99], mp1_res[100], mp1_res[110], mp1_res[111], mp1_res[112], mp1_res[123], mp1_res[125], mp1_res[127]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[51]));
    dotproduct15 operation_conv729(.clk (clk), .rst (rst), .g_input ({mp1_res[72], mp1_res[73], mp1_res[74], mp1_res[75], mp1_res[86], mp1_res[87], mp1_res[89], mp1_res[100], mp1_res[101], mp1_res[111], mp1_res[112], mp1_res[113], mp1_res[124], mp1_res[126], mp1_res[128]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[52]));
    dotproduct15 operation_conv730(.clk (clk), .rst (rst), .g_input ({mp1_res[73], mp1_res[74], mp1_res[75], mp1_res[76], mp1_res[87], mp1_res[88], mp1_res[90], mp1_res[101], mp1_res[102], mp1_res[112], mp1_res[113], mp1_res[114], mp1_res[125], mp1_res[127], mp1_res[129]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[53]));
    dotproduct15 operation_conv731(.clk (clk), .rst (rst), .g_input ({mp1_res[78], mp1_res[79], mp1_res[80], mp1_res[81], mp1_res[92], mp1_res[93], mp1_res[95], mp1_res[106], mp1_res[107], mp1_res[117], mp1_res[118], mp1_res[119], mp1_res[130], mp1_res[132], mp1_res[134]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[54]));
    dotproduct15 operation_conv732(.clk (clk), .rst (rst), .g_input ({mp1_res[79], mp1_res[80], mp1_res[81], mp1_res[82], mp1_res[93], mp1_res[94], mp1_res[96], mp1_res[107], mp1_res[108], mp1_res[118], mp1_res[119], mp1_res[120], mp1_res[131], mp1_res[133], mp1_res[135]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[55]));
    dotproduct15 operation_conv733(.clk (clk), .rst (rst), .g_input ({mp1_res[80], mp1_res[81], mp1_res[82], mp1_res[83], mp1_res[94], mp1_res[95], mp1_res[97], mp1_res[108], mp1_res[109], mp1_res[119], mp1_res[120], mp1_res[121], mp1_res[132], mp1_res[134], mp1_res[136]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[56]));
    dotproduct15 operation_conv734(.clk (clk), .rst (rst), .g_input ({mp1_res[81], mp1_res[82], mp1_res[83], mp1_res[84], mp1_res[95], mp1_res[96], mp1_res[98], mp1_res[109], mp1_res[110], mp1_res[120], mp1_res[121], mp1_res[122], mp1_res[133], mp1_res[135], mp1_res[137]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[57]));
    dotproduct15 operation_conv735(.clk (clk), .rst (rst), .g_input ({mp1_res[82], mp1_res[83], mp1_res[84], mp1_res[85], mp1_res[96], mp1_res[97], mp1_res[99], mp1_res[110], mp1_res[111], mp1_res[121], mp1_res[122], mp1_res[123], mp1_res[134], mp1_res[136], mp1_res[138]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[58]));
    dotproduct15 operation_conv736(.clk (clk), .rst (rst), .g_input ({mp1_res[83], mp1_res[84], mp1_res[85], mp1_res[86], mp1_res[97], mp1_res[98], mp1_res[100], mp1_res[111], mp1_res[112], mp1_res[122], mp1_res[123], mp1_res[124], mp1_res[135], mp1_res[137], mp1_res[139]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[59]));
    dotproduct15 operation_conv737(.clk (clk), .rst (rst), .g_input ({mp1_res[84], mp1_res[85], mp1_res[86], mp1_res[87], mp1_res[98], mp1_res[99], mp1_res[101], mp1_res[112], mp1_res[113], mp1_res[123], mp1_res[124], mp1_res[125], mp1_res[136], mp1_res[138], mp1_res[140]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[60]));
    dotproduct15 operation_conv738(.clk (clk), .rst (rst), .g_input ({mp1_res[85], mp1_res[86], mp1_res[87], mp1_res[88], mp1_res[99], mp1_res[100], mp1_res[102], mp1_res[113], mp1_res[114], mp1_res[124], mp1_res[125], mp1_res[126], mp1_res[137], mp1_res[139], mp1_res[141]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[61]));
    dotproduct15 operation_conv739(.clk (clk), .rst (rst), .g_input ({mp1_res[86], mp1_res[87], mp1_res[88], mp1_res[89], mp1_res[100], mp1_res[101], mp1_res[103], mp1_res[114], mp1_res[115], mp1_res[125], mp1_res[126], mp1_res[127], mp1_res[138], mp1_res[140], mp1_res[142]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[62]));
    dotproduct15 operation_conv740(.clk (clk), .rst (rst), .g_input ({mp1_res[91], mp1_res[92], mp1_res[93], mp1_res[94], mp1_res[105], mp1_res[106], mp1_res[108], mp1_res[119], mp1_res[120], mp1_res[130], mp1_res[131], mp1_res[132], mp1_res[143], mp1_res[145], mp1_res[147]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[63]));
    dotproduct15 operation_conv741(.clk (clk), .rst (rst), .g_input ({mp1_res[92], mp1_res[93], mp1_res[94], mp1_res[95], mp1_res[106], mp1_res[107], mp1_res[109], mp1_res[120], mp1_res[121], mp1_res[131], mp1_res[132], mp1_res[133], mp1_res[144], mp1_res[146], mp1_res[148]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[64]));
    dotproduct15 operation_conv742(.clk (clk), .rst (rst), .g_input ({mp1_res[93], mp1_res[94], mp1_res[95], mp1_res[96], mp1_res[107], mp1_res[108], mp1_res[110], mp1_res[121], mp1_res[122], mp1_res[132], mp1_res[133], mp1_res[134], mp1_res[145], mp1_res[147], mp1_res[149]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[65]));
    dotproduct15 operation_conv743(.clk (clk), .rst (rst), .g_input ({mp1_res[94], mp1_res[95], mp1_res[96], mp1_res[97], mp1_res[108], mp1_res[109], mp1_res[111], mp1_res[122], mp1_res[123], mp1_res[133], mp1_res[134], mp1_res[135], mp1_res[146], mp1_res[148], mp1_res[150]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[66]));
    dotproduct15 operation_conv744(.clk (clk), .rst (rst), .g_input ({mp1_res[95], mp1_res[96], mp1_res[97], mp1_res[98], mp1_res[109], mp1_res[110], mp1_res[112], mp1_res[123], mp1_res[124], mp1_res[134], mp1_res[135], mp1_res[136], mp1_res[147], mp1_res[149], mp1_res[151]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[67]));
    dotproduct15 operation_conv745(.clk (clk), .rst (rst), .g_input ({mp1_res[96], mp1_res[97], mp1_res[98], mp1_res[99], mp1_res[110], mp1_res[111], mp1_res[113], mp1_res[124], mp1_res[125], mp1_res[135], mp1_res[136], mp1_res[137], mp1_res[148], mp1_res[150], mp1_res[152]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[68]));
    dotproduct15 operation_conv746(.clk (clk), .rst (rst), .g_input ({mp1_res[97], mp1_res[98], mp1_res[99], mp1_res[100], mp1_res[111], mp1_res[112], mp1_res[114], mp1_res[125], mp1_res[126], mp1_res[136], mp1_res[137], mp1_res[138], mp1_res[149], mp1_res[151], mp1_res[153]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[69]));
    dotproduct15 operation_conv747(.clk (clk), .rst (rst), .g_input ({mp1_res[98], mp1_res[99], mp1_res[100], mp1_res[101], mp1_res[112], mp1_res[113], mp1_res[115], mp1_res[126], mp1_res[127], mp1_res[137], mp1_res[138], mp1_res[139], mp1_res[150], mp1_res[152], mp1_res[154]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[70]));
    dotproduct15 operation_conv748(.clk (clk), .rst (rst), .g_input ({mp1_res[99], mp1_res[100], mp1_res[101], mp1_res[102], mp1_res[113], mp1_res[114], mp1_res[116], mp1_res[127], mp1_res[128], mp1_res[138], mp1_res[139], mp1_res[140], mp1_res[151], mp1_res[153], mp1_res[155]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[71]));
    dotproduct15 operation_conv749(.clk (clk), .rst (rst), .g_input ({mp1_res[104], mp1_res[105], mp1_res[106], mp1_res[107], mp1_res[118], mp1_res[119], mp1_res[121], mp1_res[132], mp1_res[133], mp1_res[143], mp1_res[144], mp1_res[145], mp1_res[156], mp1_res[158], mp1_res[160]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[72]));
    dotproduct15 operation_conv750(.clk (clk), .rst (rst), .g_input ({mp1_res[105], mp1_res[106], mp1_res[107], mp1_res[108], mp1_res[119], mp1_res[120], mp1_res[122], mp1_res[133], mp1_res[134], mp1_res[144], mp1_res[145], mp1_res[146], mp1_res[157], mp1_res[159], mp1_res[161]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[73]));
    dotproduct15 operation_conv751(.clk (clk), .rst (rst), .g_input ({mp1_res[106], mp1_res[107], mp1_res[108], mp1_res[109], mp1_res[120], mp1_res[121], mp1_res[123], mp1_res[134], mp1_res[135], mp1_res[145], mp1_res[146], mp1_res[147], mp1_res[158], mp1_res[160], mp1_res[162]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[74]));
    dotproduct15 operation_conv752(.clk (clk), .rst (rst), .g_input ({mp1_res[107], mp1_res[108], mp1_res[109], mp1_res[110], mp1_res[121], mp1_res[122], mp1_res[124], mp1_res[135], mp1_res[136], mp1_res[146], mp1_res[147], mp1_res[148], mp1_res[159], mp1_res[161], mp1_res[163]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[75]));
    dotproduct15 operation_conv753(.clk (clk), .rst (rst), .g_input ({mp1_res[108], mp1_res[109], mp1_res[110], mp1_res[111], mp1_res[122], mp1_res[123], mp1_res[125], mp1_res[136], mp1_res[137], mp1_res[147], mp1_res[148], mp1_res[149], mp1_res[160], mp1_res[162], mp1_res[164]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[76]));
    dotproduct15 operation_conv754(.clk (clk), .rst (rst), .g_input ({mp1_res[109], mp1_res[110], mp1_res[111], mp1_res[112], mp1_res[123], mp1_res[124], mp1_res[126], mp1_res[137], mp1_res[138], mp1_res[148], mp1_res[149], mp1_res[150], mp1_res[161], mp1_res[163], mp1_res[165]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[77]));
    dotproduct15 operation_conv755(.clk (clk), .rst (rst), .g_input ({mp1_res[110], mp1_res[111], mp1_res[112], mp1_res[113], mp1_res[124], mp1_res[125], mp1_res[127], mp1_res[138], mp1_res[139], mp1_res[149], mp1_res[150], mp1_res[151], mp1_res[162], mp1_res[164], mp1_res[166]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[78]));
    dotproduct15 operation_conv756(.clk (clk), .rst (rst), .g_input ({mp1_res[111], mp1_res[112], mp1_res[113], mp1_res[114], mp1_res[125], mp1_res[126], mp1_res[128], mp1_res[139], mp1_res[140], mp1_res[150], mp1_res[151], mp1_res[152], mp1_res[163], mp1_res[165], mp1_res[167]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[79]));
    dotproduct15 operation_conv757(.clk (clk), .rst (rst), .g_input ({mp1_res[112], mp1_res[113], mp1_res[114], mp1_res[115], mp1_res[126], mp1_res[127], mp1_res[129], mp1_res[140], mp1_res[141], mp1_res[151], mp1_res[152], mp1_res[153], mp1_res[164], mp1_res[166], mp1_res[168]}), .e_input({e_input[9], e_input[10], e_input[11], e_input[12], e_input[15], e_input[16], e_input[18], e_input[21], e_input[22], e_input[24], e_input[25], e_input[26], e_input[29], e_input[31], e_input[33]}), .o (conv2_0_0[80]));
    assign conv2_res = {conv2_0_0};


    fc1 operation_fc1758(
        .clk   (clk),
        .rst   (rst),
        .g_input (conv2_res),
        .e_input (e_input[843:34]),
        .o     (fc1_res)
    );
    
    fc2 operation_fc2759(
        .clk   (clk),
        .rst   (rst),
        .g_input (fc1_res),
        .e_input (e_input[943:844]),
        .o     (fc2_res)
    );
    

assign o = fc2_res; 

endmodule
    